
module conv_20_13_20_1 ( clk, reset, s_data_in_x, s_valid_x, s_ready_x, 
        m_data_out_y, m_valid_y, m_ready_y );
  input [19:0] s_data_in_x;
  output [19:0] m_data_out_y;
  input clk, reset, s_valid_x, m_ready_y;
  output s_ready_x, m_valid_y;
  wire   conv_done, conv_pre_start, N29, \xmem_inst/N109 , \xmem_inst/N107 ,
         \xmem_inst/N106 , \xmem_inst/N105 , \xmem_inst/N103 ,
         \xmem_inst/N101 , \xmem_inst/N100 , \xmem_inst/N99 , \xmem_inst/N98 ,
         \xmem_inst/N97 , \xmem_inst/N95 , \xmem_inst/N94 , \xmem_inst/N93 ,
         \xmem_inst/N91 , \xmem_inst/mem[19][19] , \xmem_inst/mem[19][18] ,
         \xmem_inst/mem[19][17] , \xmem_inst/mem[19][16] ,
         \xmem_inst/mem[19][15] , \xmem_inst/mem[19][14] ,
         \xmem_inst/mem[19][13] , \xmem_inst/mem[19][12] ,
         \xmem_inst/mem[19][11] , \xmem_inst/mem[19][10] ,
         \xmem_inst/mem[19][9] , \xmem_inst/mem[19][8] ,
         \xmem_inst/mem[19][7] , \xmem_inst/mem[19][6] ,
         \xmem_inst/mem[19][5] , \xmem_inst/mem[19][4] ,
         \xmem_inst/mem[19][3] , \xmem_inst/mem[19][2] ,
         \xmem_inst/mem[19][1] , \xmem_inst/mem[19][0] ,
         \xmem_inst/mem[18][19] , \xmem_inst/mem[18][18] ,
         \xmem_inst/mem[18][17] , \xmem_inst/mem[18][16] ,
         \xmem_inst/mem[18][15] , \xmem_inst/mem[18][14] ,
         \xmem_inst/mem[18][13] , \xmem_inst/mem[18][12] ,
         \xmem_inst/mem[18][11] , \xmem_inst/mem[18][10] ,
         \xmem_inst/mem[18][9] , \xmem_inst/mem[18][8] ,
         \xmem_inst/mem[18][7] , \xmem_inst/mem[18][6] ,
         \xmem_inst/mem[18][5] , \xmem_inst/mem[18][4] ,
         \xmem_inst/mem[18][3] , \xmem_inst/mem[18][2] ,
         \xmem_inst/mem[18][1] , \xmem_inst/mem[18][0] ,
         \xmem_inst/mem[17][19] , \xmem_inst/mem[17][18] ,
         \xmem_inst/mem[17][17] , \xmem_inst/mem[17][16] ,
         \xmem_inst/mem[17][15] , \xmem_inst/mem[17][14] ,
         \xmem_inst/mem[17][13] , \xmem_inst/mem[17][12] ,
         \xmem_inst/mem[17][11] , \xmem_inst/mem[17][10] ,
         \xmem_inst/mem[17][9] , \xmem_inst/mem[17][8] ,
         \xmem_inst/mem[17][7] , \xmem_inst/mem[17][6] ,
         \xmem_inst/mem[17][5] , \xmem_inst/mem[17][4] ,
         \xmem_inst/mem[17][3] , \xmem_inst/mem[17][2] ,
         \xmem_inst/mem[17][1] , \xmem_inst/mem[17][0] ,
         \xmem_inst/mem[16][19] , \xmem_inst/mem[16][18] ,
         \xmem_inst/mem[16][17] , \xmem_inst/mem[16][16] ,
         \xmem_inst/mem[16][15] , \xmem_inst/mem[16][14] ,
         \xmem_inst/mem[16][13] , \xmem_inst/mem[16][12] ,
         \xmem_inst/mem[16][11] , \xmem_inst/mem[16][10] ,
         \xmem_inst/mem[16][9] , \xmem_inst/mem[16][8] ,
         \xmem_inst/mem[16][7] , \xmem_inst/mem[16][6] ,
         \xmem_inst/mem[16][5] , \xmem_inst/mem[16][4] ,
         \xmem_inst/mem[16][3] , \xmem_inst/mem[16][2] ,
         \xmem_inst/mem[16][1] , \xmem_inst/mem[16][0] ,
         \xmem_inst/mem[15][19] , \xmem_inst/mem[15][18] ,
         \xmem_inst/mem[15][17] , \xmem_inst/mem[15][16] ,
         \xmem_inst/mem[15][15] , \xmem_inst/mem[15][14] ,
         \xmem_inst/mem[15][13] , \xmem_inst/mem[15][12] ,
         \xmem_inst/mem[15][11] , \xmem_inst/mem[15][10] ,
         \xmem_inst/mem[15][9] , \xmem_inst/mem[15][8] ,
         \xmem_inst/mem[15][7] , \xmem_inst/mem[15][6] ,
         \xmem_inst/mem[15][5] , \xmem_inst/mem[15][4] ,
         \xmem_inst/mem[15][3] , \xmem_inst/mem[15][2] ,
         \xmem_inst/mem[15][1] , \xmem_inst/mem[15][0] ,
         \xmem_inst/mem[14][19] , \xmem_inst/mem[14][18] ,
         \xmem_inst/mem[14][17] , \xmem_inst/mem[14][16] ,
         \xmem_inst/mem[14][15] , \xmem_inst/mem[14][14] ,
         \xmem_inst/mem[14][13] , \xmem_inst/mem[14][12] ,
         \xmem_inst/mem[14][11] , \xmem_inst/mem[14][10] ,
         \xmem_inst/mem[14][9] , \xmem_inst/mem[14][8] ,
         \xmem_inst/mem[14][7] , \xmem_inst/mem[14][6] ,
         \xmem_inst/mem[14][5] , \xmem_inst/mem[14][4] ,
         \xmem_inst/mem[14][3] , \xmem_inst/mem[14][2] ,
         \xmem_inst/mem[14][1] , \xmem_inst/mem[14][0] ,
         \xmem_inst/mem[13][19] , \xmem_inst/mem[13][18] ,
         \xmem_inst/mem[13][17] , \xmem_inst/mem[13][16] ,
         \xmem_inst/mem[13][15] , \xmem_inst/mem[13][14] ,
         \xmem_inst/mem[13][13] , \xmem_inst/mem[13][12] ,
         \xmem_inst/mem[13][11] , \xmem_inst/mem[13][10] ,
         \xmem_inst/mem[13][9] , \xmem_inst/mem[13][8] ,
         \xmem_inst/mem[13][7] , \xmem_inst/mem[13][6] ,
         \xmem_inst/mem[13][5] , \xmem_inst/mem[13][4] ,
         \xmem_inst/mem[13][3] , \xmem_inst/mem[13][2] ,
         \xmem_inst/mem[13][1] , \xmem_inst/mem[13][0] ,
         \xmem_inst/mem[12][19] , \xmem_inst/mem[12][18] ,
         \xmem_inst/mem[12][17] , \xmem_inst/mem[12][16] ,
         \xmem_inst/mem[12][15] , \xmem_inst/mem[12][14] ,
         \xmem_inst/mem[12][13] , \xmem_inst/mem[12][12] ,
         \xmem_inst/mem[12][11] , \xmem_inst/mem[12][10] ,
         \xmem_inst/mem[12][9] , \xmem_inst/mem[12][8] ,
         \xmem_inst/mem[12][7] , \xmem_inst/mem[12][6] ,
         \xmem_inst/mem[12][5] , \xmem_inst/mem[12][4] ,
         \xmem_inst/mem[12][3] , \xmem_inst/mem[12][2] ,
         \xmem_inst/mem[12][1] , \xmem_inst/mem[12][0] ,
         \xmem_inst/mem[11][19] , \xmem_inst/mem[11][18] ,
         \xmem_inst/mem[11][17] , \xmem_inst/mem[11][16] ,
         \xmem_inst/mem[11][15] , \xmem_inst/mem[11][14] ,
         \xmem_inst/mem[11][13] , \xmem_inst/mem[11][12] ,
         \xmem_inst/mem[11][11] , \xmem_inst/mem[11][10] ,
         \xmem_inst/mem[11][9] , \xmem_inst/mem[11][8] ,
         \xmem_inst/mem[11][7] , \xmem_inst/mem[11][6] ,
         \xmem_inst/mem[11][5] , \xmem_inst/mem[11][4] ,
         \xmem_inst/mem[11][3] , \xmem_inst/mem[11][2] ,
         \xmem_inst/mem[11][1] , \xmem_inst/mem[11][0] ,
         \xmem_inst/mem[10][19] , \xmem_inst/mem[10][18] ,
         \xmem_inst/mem[10][17] , \xmem_inst/mem[10][16] ,
         \xmem_inst/mem[10][15] , \xmem_inst/mem[10][14] ,
         \xmem_inst/mem[10][13] , \xmem_inst/mem[10][12] ,
         \xmem_inst/mem[10][11] , \xmem_inst/mem[10][10] ,
         \xmem_inst/mem[10][9] , \xmem_inst/mem[10][8] ,
         \xmem_inst/mem[10][7] , \xmem_inst/mem[10][6] ,
         \xmem_inst/mem[10][5] , \xmem_inst/mem[10][4] ,
         \xmem_inst/mem[10][3] , \xmem_inst/mem[10][2] ,
         \xmem_inst/mem[10][1] , \xmem_inst/mem[10][0] ,
         \xmem_inst/mem[9][19] , \xmem_inst/mem[9][18] ,
         \xmem_inst/mem[9][17] , \xmem_inst/mem[9][16] ,
         \xmem_inst/mem[9][15] , \xmem_inst/mem[9][14] ,
         \xmem_inst/mem[9][13] , \xmem_inst/mem[9][12] ,
         \xmem_inst/mem[9][11] , \xmem_inst/mem[9][10] , \xmem_inst/mem[9][9] ,
         \xmem_inst/mem[9][8] , \xmem_inst/mem[9][7] , \xmem_inst/mem[9][6] ,
         \xmem_inst/mem[9][5] , \xmem_inst/mem[9][4] , \xmem_inst/mem[9][3] ,
         \xmem_inst/mem[9][2] , \xmem_inst/mem[9][1] , \xmem_inst/mem[9][0] ,
         \xmem_inst/mem[8][19] , \xmem_inst/mem[8][18] ,
         \xmem_inst/mem[8][17] , \xmem_inst/mem[8][16] ,
         \xmem_inst/mem[8][15] , \xmem_inst/mem[8][14] ,
         \xmem_inst/mem[8][13] , \xmem_inst/mem[8][12] ,
         \xmem_inst/mem[8][11] , \xmem_inst/mem[8][10] , \xmem_inst/mem[8][9] ,
         \xmem_inst/mem[8][8] , \xmem_inst/mem[8][7] , \xmem_inst/mem[8][6] ,
         \xmem_inst/mem[8][5] , \xmem_inst/mem[8][4] , \xmem_inst/mem[8][3] ,
         \xmem_inst/mem[8][2] , \xmem_inst/mem[8][1] , \xmem_inst/mem[8][0] ,
         \xmem_inst/mem[7][19] , \xmem_inst/mem[7][18] ,
         \xmem_inst/mem[7][17] , \xmem_inst/mem[7][16] ,
         \xmem_inst/mem[7][15] , \xmem_inst/mem[7][14] ,
         \xmem_inst/mem[7][13] , \xmem_inst/mem[7][12] ,
         \xmem_inst/mem[7][11] , \xmem_inst/mem[7][10] , \xmem_inst/mem[7][9] ,
         \xmem_inst/mem[7][8] , \xmem_inst/mem[7][7] , \xmem_inst/mem[7][6] ,
         \xmem_inst/mem[7][5] , \xmem_inst/mem[7][4] , \xmem_inst/mem[7][3] ,
         \xmem_inst/mem[7][2] , \xmem_inst/mem[7][1] , \xmem_inst/mem[7][0] ,
         \xmem_inst/mem[6][19] , \xmem_inst/mem[6][18] ,
         \xmem_inst/mem[6][17] , \xmem_inst/mem[6][16] ,
         \xmem_inst/mem[6][15] , \xmem_inst/mem[6][14] ,
         \xmem_inst/mem[6][13] , \xmem_inst/mem[6][12] ,
         \xmem_inst/mem[6][11] , \xmem_inst/mem[6][10] , \xmem_inst/mem[6][9] ,
         \xmem_inst/mem[6][8] , \xmem_inst/mem[6][7] , \xmem_inst/mem[6][6] ,
         \xmem_inst/mem[6][5] , \xmem_inst/mem[6][4] , \xmem_inst/mem[6][3] ,
         \xmem_inst/mem[6][2] , \xmem_inst/mem[6][1] , \xmem_inst/mem[6][0] ,
         \xmem_inst/mem[5][19] , \xmem_inst/mem[5][18] ,
         \xmem_inst/mem[5][17] , \xmem_inst/mem[5][16] ,
         \xmem_inst/mem[5][15] , \xmem_inst/mem[5][14] ,
         \xmem_inst/mem[5][13] , \xmem_inst/mem[5][12] ,
         \xmem_inst/mem[5][11] , \xmem_inst/mem[5][10] , \xmem_inst/mem[5][9] ,
         \xmem_inst/mem[5][8] , \xmem_inst/mem[5][7] , \xmem_inst/mem[5][6] ,
         \xmem_inst/mem[5][5] , \xmem_inst/mem[5][4] , \xmem_inst/mem[5][3] ,
         \xmem_inst/mem[5][2] , \xmem_inst/mem[5][1] , \xmem_inst/mem[5][0] ,
         \xmem_inst/mem[4][19] , \xmem_inst/mem[4][18] ,
         \xmem_inst/mem[4][17] , \xmem_inst/mem[4][16] ,
         \xmem_inst/mem[4][15] , \xmem_inst/mem[4][14] ,
         \xmem_inst/mem[4][13] , \xmem_inst/mem[4][12] ,
         \xmem_inst/mem[4][11] , \xmem_inst/mem[4][10] , \xmem_inst/mem[4][9] ,
         \xmem_inst/mem[4][8] , \xmem_inst/mem[4][7] , \xmem_inst/mem[4][6] ,
         \xmem_inst/mem[4][5] , \xmem_inst/mem[4][4] , \xmem_inst/mem[4][3] ,
         \xmem_inst/mem[4][2] , \xmem_inst/mem[4][1] , \xmem_inst/mem[4][0] ,
         \xmem_inst/mem[3][19] , \xmem_inst/mem[3][18] ,
         \xmem_inst/mem[3][17] , \xmem_inst/mem[3][16] ,
         \xmem_inst/mem[3][15] , \xmem_inst/mem[3][14] ,
         \xmem_inst/mem[3][13] , \xmem_inst/mem[3][12] ,
         \xmem_inst/mem[3][11] , \xmem_inst/mem[3][10] , \xmem_inst/mem[3][9] ,
         \xmem_inst/mem[3][8] , \xmem_inst/mem[3][7] , \xmem_inst/mem[3][6] ,
         \xmem_inst/mem[3][5] , \xmem_inst/mem[3][4] , \xmem_inst/mem[3][3] ,
         \xmem_inst/mem[3][2] , \xmem_inst/mem[3][1] , \xmem_inst/mem[3][0] ,
         \xmem_inst/mem[2][19] , \xmem_inst/mem[2][18] ,
         \xmem_inst/mem[2][17] , \xmem_inst/mem[2][16] ,
         \xmem_inst/mem[2][15] , \xmem_inst/mem[2][14] ,
         \xmem_inst/mem[2][13] , \xmem_inst/mem[2][12] ,
         \xmem_inst/mem[2][11] , \xmem_inst/mem[2][10] , \xmem_inst/mem[2][9] ,
         \xmem_inst/mem[2][8] , \xmem_inst/mem[2][7] , \xmem_inst/mem[2][6] ,
         \xmem_inst/mem[2][5] , \xmem_inst/mem[2][4] , \xmem_inst/mem[2][3] ,
         \xmem_inst/mem[2][2] , \xmem_inst/mem[2][1] , \xmem_inst/mem[2][0] ,
         \xmem_inst/mem[1][19] , \xmem_inst/mem[1][18] ,
         \xmem_inst/mem[1][17] , \xmem_inst/mem[1][16] ,
         \xmem_inst/mem[1][15] , \xmem_inst/mem[1][14] ,
         \xmem_inst/mem[1][13] , \xmem_inst/mem[1][12] ,
         \xmem_inst/mem[1][11] , \xmem_inst/mem[1][10] , \xmem_inst/mem[1][9] ,
         \xmem_inst/mem[1][8] , \xmem_inst/mem[1][7] , \xmem_inst/mem[1][6] ,
         \xmem_inst/mem[1][5] , \xmem_inst/mem[1][4] , \xmem_inst/mem[1][3] ,
         \xmem_inst/mem[1][2] , \xmem_inst/mem[1][1] , \xmem_inst/mem[1][0] ,
         \xmem_inst/mem[0][19] , \xmem_inst/mem[0][18] ,
         \xmem_inst/mem[0][17] , \xmem_inst/mem[0][16] ,
         \xmem_inst/mem[0][15] , \xmem_inst/mem[0][14] ,
         \xmem_inst/mem[0][13] , \xmem_inst/mem[0][12] ,
         \xmem_inst/mem[0][11] , \xmem_inst/mem[0][10] , \xmem_inst/mem[0][9] ,
         \xmem_inst/mem[0][8] , \xmem_inst/mem[0][7] , \xmem_inst/mem[0][6] ,
         \xmem_inst/mem[0][5] , \xmem_inst/mem[0][4] , \xmem_inst/mem[0][3] ,
         \xmem_inst/mem[0][2] , \xmem_inst/mem[0][1] , \xmem_inst/mem[0][0] ,
         \ctrl_conv_output_inst/N77 , \ctrl_conv_output_inst/N74 ,
         \ctrl_conv_output_inst/m_pre_valid_y ,
         \ctrl_conv_output_inst/conv_start_accum ,
         \ctrl_conv_output_inst/m_pre_pre_valid_y , n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, \DP_OP_485J1_122_4413/n1657 ,
         \DP_OP_485J1_122_4413/n1656 , \DP_OP_485J1_122_4413/n1655 ,
         \DP_OP_485J1_122_4413/n1204 , n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391;
  wire   [4:0] xmem_addr;
  wire   [19:0] xmem_data;
  wire   [3:0] fmem_addr;
  wire   [19:0] fmem_data;
  wire   [4:0] \ctrl_conv_output_inst/cnt_conv ;
  wire   [19:0] \mac_unit_inst/adder_reg ;
  wire   [19:0] \mac_unit_inst/x_mult_f_reg ;
  assign m_data_out_y[19] = 1'b0;

  DFF_X1 \ctrl_conv_output_inst/conv_done_reg  ( .D(
        \ctrl_conv_output_inst/N77 ), .CK(clk), .Q(conv_done) );
  DFF_X1 \fmem_addr_reg[3]  ( .D(n923), .CK(clk), .Q(fmem_addr[3]), .QN(n3339)
         );
  DFF_X1 \ctrl_conv_output_inst/m_pre_pre_valid_y_reg  ( .D(n1339), .CK(clk), 
        .Q(\ctrl_conv_output_inst/m_pre_pre_valid_y ), .QN(n3344) );
  DFF_X1 \ctrl_conv_output_inst/m_pre_valid_y_reg  ( .D(n911), .CK(clk), .Q(
        \ctrl_conv_output_inst/m_pre_valid_y ), .QN(n3336) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[4]  ( .D(n1338), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [4]), .QN(n3337) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[0]  ( .D(n1337), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [0]), .QN(n3333) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[1]  ( .D(n1336), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [1]), .QN(n3343) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[2]  ( .D(n1335), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [2]), .QN(n3341) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[3]  ( .D(n1334), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [3]), .QN(n3342) );
  DFF_X1 \ctrl_conv_output_inst/m_valid_y_reg  ( .D(n1333), .CK(clk), .Q(
        m_valid_y) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[4]  ( .D(n1327), .CK(clk), .Q(
        xmem_addr[4]), .QN(n3334) );
  DFF_X1 \ctrl_xmem_write_inst/s_ready_reg  ( .D(n1332), .CK(clk), .Q(
        s_ready_x), .QN(n3367) );
  DFF_X1 conv_pre_start_reg ( .D(N29), .CK(clk), .Q(conv_pre_start) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[0]  ( .D(n1331), .CK(clk), .Q(
        xmem_addr[0]), .QN(n3338) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[1]  ( .D(n1330), .CK(clk), .Q(
        xmem_addr[1]), .QN(n3345) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[2]  ( .D(n1329), .CK(clk), .Q(
        xmem_addr[2]), .QN(n3340) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[3]  ( .D(n1328), .CK(clk), .Q(
        xmem_addr[3]), .QN(n3335) );
  DFF_X1 \xmem_inst/mem_reg[8][0]  ( .D(n1166), .CK(clk), .Q(
        \xmem_inst/mem[8][0] ) );
  DFF_X1 \xmem_inst/mem_reg[8][1]  ( .D(n1165), .CK(clk), .Q(
        \xmem_inst/mem[8][1] ) );
  DFF_X1 \xmem_inst/mem_reg[8][2]  ( .D(n1164), .CK(clk), .Q(
        \xmem_inst/mem[8][2] ) );
  DFF_X1 \xmem_inst/mem_reg[8][3]  ( .D(n1163), .CK(clk), .Q(
        \xmem_inst/mem[8][3] ) );
  DFF_X1 \xmem_inst/mem_reg[8][4]  ( .D(n1162), .CK(clk), .Q(
        \xmem_inst/mem[8][4] ) );
  DFF_X1 \xmem_inst/mem_reg[8][5]  ( .D(n1161), .CK(clk), .Q(
        \xmem_inst/mem[8][5] ) );
  DFF_X1 \xmem_inst/mem_reg[8][6]  ( .D(n1160), .CK(clk), .Q(
        \xmem_inst/mem[8][6] ) );
  DFF_X1 \xmem_inst/mem_reg[8][7]  ( .D(n1159), .CK(clk), .Q(
        \xmem_inst/mem[8][7] ) );
  DFF_X1 \xmem_inst/mem_reg[8][8]  ( .D(n1158), .CK(clk), .Q(
        \xmem_inst/mem[8][8] ) );
  DFF_X1 \xmem_inst/mem_reg[8][9]  ( .D(n1157), .CK(clk), .Q(
        \xmem_inst/mem[8][9] ) );
  DFF_X1 \xmem_inst/mem_reg[8][10]  ( .D(n1156), .CK(clk), .Q(
        \xmem_inst/mem[8][10] ) );
  DFF_X1 \xmem_inst/mem_reg[8][11]  ( .D(n1155), .CK(clk), .Q(
        \xmem_inst/mem[8][11] ) );
  DFF_X1 \xmem_inst/mem_reg[8][12]  ( .D(n1154), .CK(clk), .Q(
        \xmem_inst/mem[8][12] ) );
  DFF_X1 \xmem_inst/mem_reg[8][13]  ( .D(n1153), .CK(clk), .Q(
        \xmem_inst/mem[8][13] ) );
  DFF_X1 \xmem_inst/mem_reg[8][14]  ( .D(n1152), .CK(clk), .Q(
        \xmem_inst/mem[8][14] ) );
  DFF_X1 \xmem_inst/mem_reg[8][15]  ( .D(n1151), .CK(clk), .Q(
        \xmem_inst/mem[8][15] ) );
  DFF_X1 \xmem_inst/mem_reg[8][16]  ( .D(n1150), .CK(clk), .Q(
        \xmem_inst/mem[8][16] ) );
  DFF_X1 \xmem_inst/mem_reg[8][17]  ( .D(n1149), .CK(clk), .Q(
        \xmem_inst/mem[8][17] ) );
  DFF_X1 \xmem_inst/mem_reg[8][18]  ( .D(n1148), .CK(clk), .Q(
        \xmem_inst/mem[8][18] ) );
  DFF_X1 \xmem_inst/mem_reg[8][19]  ( .D(n1147), .CK(clk), .Q(
        \xmem_inst/mem[8][19] ) );
  DFF_X1 \xmem_inst/mem_reg[9][0]  ( .D(n1146), .CK(clk), .Q(
        \xmem_inst/mem[9][0] ) );
  DFF_X1 \xmem_inst/mem_reg[9][1]  ( .D(n1145), .CK(clk), .Q(
        \xmem_inst/mem[9][1] ) );
  DFF_X1 \xmem_inst/mem_reg[9][2]  ( .D(n1144), .CK(clk), .Q(
        \xmem_inst/mem[9][2] ) );
  DFF_X1 \xmem_inst/mem_reg[9][3]  ( .D(n1143), .CK(clk), .Q(
        \xmem_inst/mem[9][3] ) );
  DFF_X1 \xmem_inst/mem_reg[9][4]  ( .D(n1142), .CK(clk), .Q(
        \xmem_inst/mem[9][4] ) );
  DFF_X1 \xmem_inst/mem_reg[9][5]  ( .D(n1141), .CK(clk), .Q(
        \xmem_inst/mem[9][5] ) );
  DFF_X1 \xmem_inst/mem_reg[9][6]  ( .D(n1140), .CK(clk), .Q(
        \xmem_inst/mem[9][6] ) );
  DFF_X1 \xmem_inst/mem_reg[9][7]  ( .D(n1139), .CK(clk), .Q(
        \xmem_inst/mem[9][7] ) );
  DFF_X1 \xmem_inst/mem_reg[9][8]  ( .D(n1138), .CK(clk), .Q(
        \xmem_inst/mem[9][8] ) );
  DFF_X1 \xmem_inst/mem_reg[9][9]  ( .D(n1137), .CK(clk), .Q(
        \xmem_inst/mem[9][9] ) );
  DFF_X1 \xmem_inst/mem_reg[9][10]  ( .D(n1136), .CK(clk), .Q(
        \xmem_inst/mem[9][10] ) );
  DFF_X1 \xmem_inst/mem_reg[9][11]  ( .D(n1135), .CK(clk), .Q(
        \xmem_inst/mem[9][11] ) );
  DFF_X1 \xmem_inst/mem_reg[9][12]  ( .D(n1134), .CK(clk), .Q(
        \xmem_inst/mem[9][12] ) );
  DFF_X1 \xmem_inst/mem_reg[9][13]  ( .D(n1133), .CK(clk), .Q(
        \xmem_inst/mem[9][13] ) );
  DFF_X1 \xmem_inst/mem_reg[9][14]  ( .D(n1132), .CK(clk), .Q(
        \xmem_inst/mem[9][14] ) );
  DFF_X1 \xmem_inst/mem_reg[9][15]  ( .D(n1131), .CK(clk), .Q(
        \xmem_inst/mem[9][15] ) );
  DFF_X1 \xmem_inst/mem_reg[9][16]  ( .D(n1130), .CK(clk), .Q(
        \xmem_inst/mem[9][16] ) );
  DFF_X1 \xmem_inst/mem_reg[9][17]  ( .D(n1129), .CK(clk), .Q(
        \xmem_inst/mem[9][17] ) );
  DFF_X1 \xmem_inst/mem_reg[9][18]  ( .D(n1128), .CK(clk), .Q(
        \xmem_inst/mem[9][18] ) );
  DFF_X1 \xmem_inst/mem_reg[9][19]  ( .D(n1127), .CK(clk), .Q(
        \xmem_inst/mem[9][19] ) );
  DFF_X1 \xmem_inst/mem_reg[10][0]  ( .D(n1126), .CK(clk), .Q(
        \xmem_inst/mem[10][0] ) );
  DFF_X1 \xmem_inst/mem_reg[10][1]  ( .D(n1125), .CK(clk), .Q(
        \xmem_inst/mem[10][1] ) );
  DFF_X1 \xmem_inst/mem_reg[10][2]  ( .D(n1124), .CK(clk), .Q(
        \xmem_inst/mem[10][2] ) );
  DFF_X1 \xmem_inst/mem_reg[10][3]  ( .D(n1123), .CK(clk), .Q(
        \xmem_inst/mem[10][3] ) );
  DFF_X1 \xmem_inst/mem_reg[10][4]  ( .D(n1122), .CK(clk), .Q(
        \xmem_inst/mem[10][4] ) );
  DFF_X1 \xmem_inst/mem_reg[10][5]  ( .D(n1121), .CK(clk), .Q(
        \xmem_inst/mem[10][5] ) );
  DFF_X1 \xmem_inst/mem_reg[10][6]  ( .D(n1120), .CK(clk), .Q(
        \xmem_inst/mem[10][6] ) );
  DFF_X1 \xmem_inst/mem_reg[10][7]  ( .D(n1119), .CK(clk), .Q(
        \xmem_inst/mem[10][7] ) );
  DFF_X1 \xmem_inst/mem_reg[10][8]  ( .D(n1118), .CK(clk), .Q(
        \xmem_inst/mem[10][8] ) );
  DFF_X1 \xmem_inst/mem_reg[10][9]  ( .D(n1117), .CK(clk), .Q(
        \xmem_inst/mem[10][9] ) );
  DFF_X1 \xmem_inst/mem_reg[10][10]  ( .D(n1116), .CK(clk), .Q(
        \xmem_inst/mem[10][10] ) );
  DFF_X1 \xmem_inst/mem_reg[10][11]  ( .D(n1115), .CK(clk), .Q(
        \xmem_inst/mem[10][11] ) );
  DFF_X1 \xmem_inst/mem_reg[10][12]  ( .D(n1114), .CK(clk), .Q(
        \xmem_inst/mem[10][12] ) );
  DFF_X1 \xmem_inst/mem_reg[10][13]  ( .D(n1113), .CK(clk), .Q(
        \xmem_inst/mem[10][13] ) );
  DFF_X1 \xmem_inst/mem_reg[10][14]  ( .D(n1112), .CK(clk), .Q(
        \xmem_inst/mem[10][14] ) );
  DFF_X1 \xmem_inst/mem_reg[10][15]  ( .D(n1111), .CK(clk), .Q(
        \xmem_inst/mem[10][15] ) );
  DFF_X1 \xmem_inst/mem_reg[10][16]  ( .D(n1110), .CK(clk), .Q(
        \xmem_inst/mem[10][16] ) );
  DFF_X1 \xmem_inst/mem_reg[10][17]  ( .D(n1109), .CK(clk), .Q(
        \xmem_inst/mem[10][17] ) );
  DFF_X1 \xmem_inst/mem_reg[10][18]  ( .D(n1108), .CK(clk), .Q(
        \xmem_inst/mem[10][18] ) );
  DFF_X1 \xmem_inst/mem_reg[10][19]  ( .D(n1107), .CK(clk), .Q(
        \xmem_inst/mem[10][19] ) );
  DFF_X1 \xmem_inst/mem_reg[11][0]  ( .D(n1106), .CK(clk), .Q(
        \xmem_inst/mem[11][0] ) );
  DFF_X1 \xmem_inst/mem_reg[11][1]  ( .D(n1105), .CK(clk), .Q(
        \xmem_inst/mem[11][1] ) );
  DFF_X1 \xmem_inst/mem_reg[11][2]  ( .D(n1104), .CK(clk), .Q(
        \xmem_inst/mem[11][2] ) );
  DFF_X1 \xmem_inst/mem_reg[11][3]  ( .D(n1103), .CK(clk), .Q(
        \xmem_inst/mem[11][3] ) );
  DFF_X1 \xmem_inst/mem_reg[11][4]  ( .D(n1102), .CK(clk), .Q(
        \xmem_inst/mem[11][4] ) );
  DFF_X1 \xmem_inst/mem_reg[11][5]  ( .D(n1101), .CK(clk), .Q(
        \xmem_inst/mem[11][5] ) );
  DFF_X1 \xmem_inst/mem_reg[11][6]  ( .D(n1100), .CK(clk), .Q(
        \xmem_inst/mem[11][6] ) );
  DFF_X1 \xmem_inst/mem_reg[11][7]  ( .D(n1099), .CK(clk), .Q(
        \xmem_inst/mem[11][7] ) );
  DFF_X1 \xmem_inst/mem_reg[11][8]  ( .D(n1098), .CK(clk), .Q(
        \xmem_inst/mem[11][8] ) );
  DFF_X1 \xmem_inst/mem_reg[11][9]  ( .D(n1097), .CK(clk), .Q(
        \xmem_inst/mem[11][9] ) );
  DFF_X1 \xmem_inst/mem_reg[11][10]  ( .D(n1096), .CK(clk), .Q(
        \xmem_inst/mem[11][10] ) );
  DFF_X1 \xmem_inst/mem_reg[11][11]  ( .D(n1095), .CK(clk), .Q(
        \xmem_inst/mem[11][11] ) );
  DFF_X1 \xmem_inst/mem_reg[11][12]  ( .D(n1094), .CK(clk), .Q(
        \xmem_inst/mem[11][12] ) );
  DFF_X1 \xmem_inst/mem_reg[11][13]  ( .D(n1093), .CK(clk), .Q(
        \xmem_inst/mem[11][13] ) );
  DFF_X1 \xmem_inst/mem_reg[11][14]  ( .D(n1092), .CK(clk), .Q(
        \xmem_inst/mem[11][14] ) );
  DFF_X1 \xmem_inst/mem_reg[11][15]  ( .D(n1091), .CK(clk), .Q(
        \xmem_inst/mem[11][15] ) );
  DFF_X1 \xmem_inst/mem_reg[11][16]  ( .D(n1090), .CK(clk), .Q(
        \xmem_inst/mem[11][16] ) );
  DFF_X1 \xmem_inst/mem_reg[11][17]  ( .D(n1089), .CK(clk), .Q(
        \xmem_inst/mem[11][17] ) );
  DFF_X1 \xmem_inst/mem_reg[11][18]  ( .D(n1088), .CK(clk), .Q(
        \xmem_inst/mem[11][18] ) );
  DFF_X1 \xmem_inst/mem_reg[11][19]  ( .D(n1087), .CK(clk), .Q(
        \xmem_inst/mem[11][19] ) );
  DFF_X1 \xmem_inst/mem_reg[12][0]  ( .D(n1086), .CK(clk), .Q(
        \xmem_inst/mem[12][0] ) );
  DFF_X1 \xmem_inst/mem_reg[12][1]  ( .D(n1085), .CK(clk), .Q(
        \xmem_inst/mem[12][1] ) );
  DFF_X1 \xmem_inst/mem_reg[12][2]  ( .D(n1084), .CK(clk), .Q(
        \xmem_inst/mem[12][2] ) );
  DFF_X1 \xmem_inst/mem_reg[12][3]  ( .D(n1083), .CK(clk), .Q(
        \xmem_inst/mem[12][3] ) );
  DFF_X1 \xmem_inst/mem_reg[12][4]  ( .D(n1082), .CK(clk), .Q(
        \xmem_inst/mem[12][4] ) );
  DFF_X1 \xmem_inst/mem_reg[12][5]  ( .D(n1081), .CK(clk), .Q(
        \xmem_inst/mem[12][5] ) );
  DFF_X1 \xmem_inst/mem_reg[12][6]  ( .D(n1080), .CK(clk), .Q(
        \xmem_inst/mem[12][6] ) );
  DFF_X1 \xmem_inst/mem_reg[12][7]  ( .D(n1079), .CK(clk), .Q(
        \xmem_inst/mem[12][7] ) );
  DFF_X1 \xmem_inst/mem_reg[12][8]  ( .D(n1078), .CK(clk), .Q(
        \xmem_inst/mem[12][8] ) );
  DFF_X1 \xmem_inst/mem_reg[12][9]  ( .D(n1077), .CK(clk), .Q(
        \xmem_inst/mem[12][9] ) );
  DFF_X1 \xmem_inst/mem_reg[12][10]  ( .D(n1076), .CK(clk), .Q(
        \xmem_inst/mem[12][10] ) );
  DFF_X1 \xmem_inst/mem_reg[12][11]  ( .D(n1075), .CK(clk), .Q(
        \xmem_inst/mem[12][11] ) );
  DFF_X1 \xmem_inst/mem_reg[12][12]  ( .D(n1074), .CK(clk), .Q(
        \xmem_inst/mem[12][12] ) );
  DFF_X1 \xmem_inst/mem_reg[12][13]  ( .D(n1073), .CK(clk), .Q(
        \xmem_inst/mem[12][13] ) );
  DFF_X1 \xmem_inst/mem_reg[12][14]  ( .D(n1072), .CK(clk), .Q(
        \xmem_inst/mem[12][14] ) );
  DFF_X1 \xmem_inst/mem_reg[12][15]  ( .D(n1071), .CK(clk), .Q(
        \xmem_inst/mem[12][15] ) );
  DFF_X1 \xmem_inst/mem_reg[12][16]  ( .D(n1070), .CK(clk), .Q(
        \xmem_inst/mem[12][16] ) );
  DFF_X1 \xmem_inst/mem_reg[12][17]  ( .D(n1069), .CK(clk), .Q(
        \xmem_inst/mem[12][17] ) );
  DFF_X1 \xmem_inst/mem_reg[12][18]  ( .D(n1068), .CK(clk), .Q(
        \xmem_inst/mem[12][18] ) );
  DFF_X1 \xmem_inst/mem_reg[12][19]  ( .D(n1067), .CK(clk), .Q(
        \xmem_inst/mem[12][19] ) );
  DFF_X1 \xmem_inst/mem_reg[13][0]  ( .D(n1066), .CK(clk), .Q(
        \xmem_inst/mem[13][0] ) );
  DFF_X1 \xmem_inst/mem_reg[13][1]  ( .D(n1065), .CK(clk), .Q(
        \xmem_inst/mem[13][1] ) );
  DFF_X1 \xmem_inst/mem_reg[13][2]  ( .D(n1064), .CK(clk), .Q(
        \xmem_inst/mem[13][2] ) );
  DFF_X1 \xmem_inst/mem_reg[13][3]  ( .D(n1063), .CK(clk), .Q(
        \xmem_inst/mem[13][3] ) );
  DFF_X1 \xmem_inst/mem_reg[13][4]  ( .D(n1062), .CK(clk), .Q(
        \xmem_inst/mem[13][4] ) );
  DFF_X1 \xmem_inst/mem_reg[13][5]  ( .D(n1061), .CK(clk), .Q(
        \xmem_inst/mem[13][5] ) );
  DFF_X1 \xmem_inst/mem_reg[13][6]  ( .D(n1060), .CK(clk), .Q(
        \xmem_inst/mem[13][6] ) );
  DFF_X1 \xmem_inst/mem_reg[13][7]  ( .D(n1059), .CK(clk), .Q(
        \xmem_inst/mem[13][7] ) );
  DFF_X1 \xmem_inst/mem_reg[13][8]  ( .D(n1058), .CK(clk), .Q(
        \xmem_inst/mem[13][8] ) );
  DFF_X1 \xmem_inst/mem_reg[13][9]  ( .D(n1057), .CK(clk), .Q(
        \xmem_inst/mem[13][9] ) );
  DFF_X1 \xmem_inst/mem_reg[13][10]  ( .D(n1056), .CK(clk), .Q(
        \xmem_inst/mem[13][10] ) );
  DFF_X1 \xmem_inst/mem_reg[13][11]  ( .D(n1055), .CK(clk), .Q(
        \xmem_inst/mem[13][11] ) );
  DFF_X1 \xmem_inst/mem_reg[13][12]  ( .D(n1054), .CK(clk), .Q(
        \xmem_inst/mem[13][12] ) );
  DFF_X1 \xmem_inst/mem_reg[13][13]  ( .D(n1053), .CK(clk), .Q(
        \xmem_inst/mem[13][13] ) );
  DFF_X1 \xmem_inst/mem_reg[13][14]  ( .D(n1052), .CK(clk), .Q(
        \xmem_inst/mem[13][14] ) );
  DFF_X1 \xmem_inst/mem_reg[13][15]  ( .D(n1051), .CK(clk), .Q(
        \xmem_inst/mem[13][15] ) );
  DFF_X1 \xmem_inst/mem_reg[13][16]  ( .D(n1050), .CK(clk), .Q(
        \xmem_inst/mem[13][16] ) );
  DFF_X1 \xmem_inst/mem_reg[13][17]  ( .D(n1049), .CK(clk), .Q(
        \xmem_inst/mem[13][17] ) );
  DFF_X1 \xmem_inst/mem_reg[13][18]  ( .D(n1048), .CK(clk), .Q(
        \xmem_inst/mem[13][18] ) );
  DFF_X1 \xmem_inst/mem_reg[13][19]  ( .D(n1047), .CK(clk), .Q(
        \xmem_inst/mem[13][19] ) );
  DFF_X1 \xmem_inst/mem_reg[14][0]  ( .D(n1046), .CK(clk), .Q(
        \xmem_inst/mem[14][0] ) );
  DFF_X1 \xmem_inst/mem_reg[14][1]  ( .D(n1045), .CK(clk), .Q(
        \xmem_inst/mem[14][1] ) );
  DFF_X1 \xmem_inst/mem_reg[14][2]  ( .D(n1044), .CK(clk), .Q(
        \xmem_inst/mem[14][2] ) );
  DFF_X1 \xmem_inst/mem_reg[14][3]  ( .D(n1043), .CK(clk), .Q(
        \xmem_inst/mem[14][3] ) );
  DFF_X1 \xmem_inst/mem_reg[14][4]  ( .D(n1042), .CK(clk), .Q(
        \xmem_inst/mem[14][4] ) );
  DFF_X1 \xmem_inst/mem_reg[14][5]  ( .D(n1041), .CK(clk), .Q(
        \xmem_inst/mem[14][5] ) );
  DFF_X1 \xmem_inst/mem_reg[14][6]  ( .D(n1040), .CK(clk), .Q(
        \xmem_inst/mem[14][6] ) );
  DFF_X1 \xmem_inst/mem_reg[14][7]  ( .D(n1039), .CK(clk), .Q(
        \xmem_inst/mem[14][7] ) );
  DFF_X1 \xmem_inst/mem_reg[14][8]  ( .D(n1038), .CK(clk), .Q(
        \xmem_inst/mem[14][8] ) );
  DFF_X1 \xmem_inst/mem_reg[14][9]  ( .D(n1037), .CK(clk), .Q(
        \xmem_inst/mem[14][9] ) );
  DFF_X1 \xmem_inst/mem_reg[14][10]  ( .D(n1036), .CK(clk), .Q(
        \xmem_inst/mem[14][10] ) );
  DFF_X1 \xmem_inst/mem_reg[14][11]  ( .D(n1035), .CK(clk), .Q(
        \xmem_inst/mem[14][11] ) );
  DFF_X1 \xmem_inst/mem_reg[14][12]  ( .D(n1034), .CK(clk), .Q(
        \xmem_inst/mem[14][12] ) );
  DFF_X1 \xmem_inst/mem_reg[14][13]  ( .D(n1033), .CK(clk), .Q(
        \xmem_inst/mem[14][13] ) );
  DFF_X1 \xmem_inst/mem_reg[14][14]  ( .D(n1032), .CK(clk), .Q(
        \xmem_inst/mem[14][14] ) );
  DFF_X1 \xmem_inst/mem_reg[14][15]  ( .D(n1031), .CK(clk), .Q(
        \xmem_inst/mem[14][15] ) );
  DFF_X1 \xmem_inst/mem_reg[14][16]  ( .D(n1030), .CK(clk), .Q(
        \xmem_inst/mem[14][16] ) );
  DFF_X1 \xmem_inst/mem_reg[14][17]  ( .D(n1029), .CK(clk), .Q(
        \xmem_inst/mem[14][17] ) );
  DFF_X1 \xmem_inst/mem_reg[14][18]  ( .D(n1028), .CK(clk), .Q(
        \xmem_inst/mem[14][18] ) );
  DFF_X1 \xmem_inst/mem_reg[14][19]  ( .D(n1027), .CK(clk), .Q(
        \xmem_inst/mem[14][19] ) );
  DFF_X1 \xmem_inst/mem_reg[15][0]  ( .D(n1026), .CK(clk), .Q(
        \xmem_inst/mem[15][0] ) );
  DFF_X1 \xmem_inst/mem_reg[15][1]  ( .D(n1025), .CK(clk), .Q(
        \xmem_inst/mem[15][1] ) );
  DFF_X1 \xmem_inst/mem_reg[15][2]  ( .D(n1024), .CK(clk), .Q(
        \xmem_inst/mem[15][2] ) );
  DFF_X1 \xmem_inst/mem_reg[15][3]  ( .D(n1023), .CK(clk), .Q(
        \xmem_inst/mem[15][3] ) );
  DFF_X1 \xmem_inst/mem_reg[15][4]  ( .D(n1022), .CK(clk), .Q(
        \xmem_inst/mem[15][4] ) );
  DFF_X1 \xmem_inst/mem_reg[15][5]  ( .D(n1021), .CK(clk), .Q(
        \xmem_inst/mem[15][5] ) );
  DFF_X1 \xmem_inst/mem_reg[15][6]  ( .D(n1020), .CK(clk), .Q(
        \xmem_inst/mem[15][6] ) );
  DFF_X1 \xmem_inst/mem_reg[15][7]  ( .D(n1019), .CK(clk), .Q(
        \xmem_inst/mem[15][7] ) );
  DFF_X1 \xmem_inst/mem_reg[15][8]  ( .D(n1018), .CK(clk), .Q(
        \xmem_inst/mem[15][8] ) );
  DFF_X1 \xmem_inst/mem_reg[15][9]  ( .D(n1017), .CK(clk), .Q(
        \xmem_inst/mem[15][9] ) );
  DFF_X1 \xmem_inst/mem_reg[15][10]  ( .D(n1016), .CK(clk), .Q(
        \xmem_inst/mem[15][10] ) );
  DFF_X1 \xmem_inst/mem_reg[15][11]  ( .D(n1015), .CK(clk), .Q(
        \xmem_inst/mem[15][11] ) );
  DFF_X1 \xmem_inst/mem_reg[15][12]  ( .D(n1014), .CK(clk), .Q(
        \xmem_inst/mem[15][12] ) );
  DFF_X1 \xmem_inst/mem_reg[15][13]  ( .D(n1013), .CK(clk), .Q(
        \xmem_inst/mem[15][13] ) );
  DFF_X1 \xmem_inst/mem_reg[15][14]  ( .D(n1012), .CK(clk), .Q(
        \xmem_inst/mem[15][14] ) );
  DFF_X1 \xmem_inst/mem_reg[15][15]  ( .D(n1011), .CK(clk), .Q(
        \xmem_inst/mem[15][15] ) );
  DFF_X1 \xmem_inst/mem_reg[15][16]  ( .D(n1010), .CK(clk), .Q(
        \xmem_inst/mem[15][16] ) );
  DFF_X1 \xmem_inst/mem_reg[15][17]  ( .D(n1009), .CK(clk), .Q(
        \xmem_inst/mem[15][17] ) );
  DFF_X1 \xmem_inst/mem_reg[15][18]  ( .D(n1008), .CK(clk), .Q(
        \xmem_inst/mem[15][18] ) );
  DFF_X1 \xmem_inst/mem_reg[15][19]  ( .D(n1007), .CK(clk), .Q(
        \xmem_inst/mem[15][19] ) );
  DFF_X1 \xmem_inst/mem_reg[0][0]  ( .D(n1326), .CK(clk), .Q(
        \xmem_inst/mem[0][0] ) );
  DFF_X1 \xmem_inst/mem_reg[0][1]  ( .D(n1325), .CK(clk), .Q(
        \xmem_inst/mem[0][1] ) );
  DFF_X1 \xmem_inst/mem_reg[0][2]  ( .D(n1324), .CK(clk), .Q(
        \xmem_inst/mem[0][2] ) );
  DFF_X1 \xmem_inst/mem_reg[0][3]  ( .D(n1323), .CK(clk), .Q(
        \xmem_inst/mem[0][3] ) );
  DFF_X1 \xmem_inst/mem_reg[0][4]  ( .D(n1322), .CK(clk), .Q(
        \xmem_inst/mem[0][4] ) );
  DFF_X1 \xmem_inst/mem_reg[0][5]  ( .D(n1321), .CK(clk), .Q(
        \xmem_inst/mem[0][5] ) );
  DFF_X1 \xmem_inst/mem_reg[0][6]  ( .D(n1320), .CK(clk), .Q(
        \xmem_inst/mem[0][6] ) );
  DFF_X1 \xmem_inst/mem_reg[0][7]  ( .D(n1319), .CK(clk), .Q(
        \xmem_inst/mem[0][7] ) );
  DFF_X1 \xmem_inst/mem_reg[0][8]  ( .D(n1318), .CK(clk), .Q(
        \xmem_inst/mem[0][8] ) );
  DFF_X1 \xmem_inst/mem_reg[0][9]  ( .D(n1317), .CK(clk), .Q(
        \xmem_inst/mem[0][9] ) );
  DFF_X1 \xmem_inst/mem_reg[0][10]  ( .D(n1316), .CK(clk), .Q(
        \xmem_inst/mem[0][10] ) );
  DFF_X1 \xmem_inst/mem_reg[0][11]  ( .D(n1315), .CK(clk), .Q(
        \xmem_inst/mem[0][11] ) );
  DFF_X1 \xmem_inst/mem_reg[0][12]  ( .D(n1314), .CK(clk), .Q(
        \xmem_inst/mem[0][12] ) );
  DFF_X1 \xmem_inst/mem_reg[0][13]  ( .D(n1313), .CK(clk), .Q(
        \xmem_inst/mem[0][13] ) );
  DFF_X1 \xmem_inst/mem_reg[0][14]  ( .D(n1312), .CK(clk), .Q(
        \xmem_inst/mem[0][14] ) );
  DFF_X1 \xmem_inst/mem_reg[0][15]  ( .D(n1311), .CK(clk), .Q(
        \xmem_inst/mem[0][15] ) );
  DFF_X1 \xmem_inst/mem_reg[0][16]  ( .D(n1310), .CK(clk), .Q(
        \xmem_inst/mem[0][16] ) );
  DFF_X1 \xmem_inst/mem_reg[0][17]  ( .D(n1309), .CK(clk), .Q(
        \xmem_inst/mem[0][17] ) );
  DFF_X1 \xmem_inst/mem_reg[0][18]  ( .D(n1308), .CK(clk), .Q(
        \xmem_inst/mem[0][18] ) );
  DFF_X1 \xmem_inst/mem_reg[0][19]  ( .D(n1307), .CK(clk), .Q(
        \xmem_inst/mem[0][19] ) );
  DFF_X1 \xmem_inst/mem_reg[1][0]  ( .D(n1306), .CK(clk), .Q(
        \xmem_inst/mem[1][0] ) );
  DFF_X1 \xmem_inst/mem_reg[1][1]  ( .D(n1305), .CK(clk), .Q(
        \xmem_inst/mem[1][1] ) );
  DFF_X1 \xmem_inst/mem_reg[1][2]  ( .D(n1304), .CK(clk), .Q(
        \xmem_inst/mem[1][2] ) );
  DFF_X1 \xmem_inst/mem_reg[1][3]  ( .D(n1303), .CK(clk), .Q(
        \xmem_inst/mem[1][3] ) );
  DFF_X1 \xmem_inst/mem_reg[1][4]  ( .D(n1302), .CK(clk), .Q(
        \xmem_inst/mem[1][4] ) );
  DFF_X1 \xmem_inst/mem_reg[1][5]  ( .D(n1301), .CK(clk), .Q(
        \xmem_inst/mem[1][5] ) );
  DFF_X1 \xmem_inst/mem_reg[1][6]  ( .D(n1300), .CK(clk), .Q(
        \xmem_inst/mem[1][6] ) );
  DFF_X1 \xmem_inst/mem_reg[1][7]  ( .D(n1299), .CK(clk), .Q(
        \xmem_inst/mem[1][7] ) );
  DFF_X1 \xmem_inst/mem_reg[1][8]  ( .D(n1298), .CK(clk), .Q(
        \xmem_inst/mem[1][8] ) );
  DFF_X1 \xmem_inst/mem_reg[1][9]  ( .D(n1297), .CK(clk), .Q(
        \xmem_inst/mem[1][9] ) );
  DFF_X1 \xmem_inst/mem_reg[1][10]  ( .D(n1296), .CK(clk), .Q(
        \xmem_inst/mem[1][10] ) );
  DFF_X1 \xmem_inst/mem_reg[1][11]  ( .D(n1295), .CK(clk), .Q(
        \xmem_inst/mem[1][11] ) );
  DFF_X1 \xmem_inst/mem_reg[1][12]  ( .D(n1294), .CK(clk), .Q(
        \xmem_inst/mem[1][12] ) );
  DFF_X1 \xmem_inst/mem_reg[1][13]  ( .D(n1293), .CK(clk), .Q(
        \xmem_inst/mem[1][13] ) );
  DFF_X1 \xmem_inst/mem_reg[1][14]  ( .D(n1292), .CK(clk), .Q(
        \xmem_inst/mem[1][14] ) );
  DFF_X1 \xmem_inst/mem_reg[1][15]  ( .D(n1291), .CK(clk), .Q(
        \xmem_inst/mem[1][15] ) );
  DFF_X1 \xmem_inst/mem_reg[1][16]  ( .D(n1290), .CK(clk), .Q(
        \xmem_inst/mem[1][16] ) );
  DFF_X1 \xmem_inst/mem_reg[1][17]  ( .D(n1289), .CK(clk), .Q(
        \xmem_inst/mem[1][17] ) );
  DFF_X1 \xmem_inst/mem_reg[1][18]  ( .D(n1288), .CK(clk), .Q(
        \xmem_inst/mem[1][18] ) );
  DFF_X1 \xmem_inst/mem_reg[1][19]  ( .D(n1287), .CK(clk), .Q(
        \xmem_inst/mem[1][19] ) );
  DFF_X1 \xmem_inst/mem_reg[2][0]  ( .D(n1286), .CK(clk), .Q(
        \xmem_inst/mem[2][0] ) );
  DFF_X1 \xmem_inst/mem_reg[2][1]  ( .D(n1285), .CK(clk), .Q(
        \xmem_inst/mem[2][1] ) );
  DFF_X1 \xmem_inst/mem_reg[2][2]  ( .D(n1284), .CK(clk), .Q(
        \xmem_inst/mem[2][2] ) );
  DFF_X1 \xmem_inst/mem_reg[2][3]  ( .D(n1283), .CK(clk), .Q(
        \xmem_inst/mem[2][3] ) );
  DFF_X1 \xmem_inst/mem_reg[2][4]  ( .D(n1282), .CK(clk), .Q(
        \xmem_inst/mem[2][4] ) );
  DFF_X1 \xmem_inst/mem_reg[2][5]  ( .D(n1281), .CK(clk), .Q(
        \xmem_inst/mem[2][5] ) );
  DFF_X1 \xmem_inst/mem_reg[2][6]  ( .D(n1280), .CK(clk), .Q(
        \xmem_inst/mem[2][6] ) );
  DFF_X1 \xmem_inst/mem_reg[2][7]  ( .D(n1279), .CK(clk), .Q(
        \xmem_inst/mem[2][7] ) );
  DFF_X1 \xmem_inst/mem_reg[2][8]  ( .D(n1278), .CK(clk), .Q(
        \xmem_inst/mem[2][8] ) );
  DFF_X1 \xmem_inst/mem_reg[2][9]  ( .D(n1277), .CK(clk), .Q(
        \xmem_inst/mem[2][9] ) );
  DFF_X1 \xmem_inst/mem_reg[2][10]  ( .D(n1276), .CK(clk), .Q(
        \xmem_inst/mem[2][10] ) );
  DFF_X1 \xmem_inst/mem_reg[2][11]  ( .D(n1275), .CK(clk), .Q(
        \xmem_inst/mem[2][11] ) );
  DFF_X1 \xmem_inst/mem_reg[2][12]  ( .D(n1274), .CK(clk), .Q(
        \xmem_inst/mem[2][12] ) );
  DFF_X1 \xmem_inst/mem_reg[2][13]  ( .D(n1273), .CK(clk), .Q(
        \xmem_inst/mem[2][13] ) );
  DFF_X1 \xmem_inst/mem_reg[2][14]  ( .D(n1272), .CK(clk), .Q(
        \xmem_inst/mem[2][14] ) );
  DFF_X1 \xmem_inst/mem_reg[2][15]  ( .D(n1271), .CK(clk), .Q(
        \xmem_inst/mem[2][15] ) );
  DFF_X1 \xmem_inst/mem_reg[2][16]  ( .D(n1270), .CK(clk), .Q(
        \xmem_inst/mem[2][16] ) );
  DFF_X1 \xmem_inst/mem_reg[2][17]  ( .D(n1269), .CK(clk), .Q(
        \xmem_inst/mem[2][17] ) );
  DFF_X1 \xmem_inst/mem_reg[2][18]  ( .D(n1268), .CK(clk), .Q(
        \xmem_inst/mem[2][18] ) );
  DFF_X1 \xmem_inst/mem_reg[2][19]  ( .D(n1267), .CK(clk), .Q(
        \xmem_inst/mem[2][19] ) );
  DFF_X1 \xmem_inst/mem_reg[3][0]  ( .D(n1266), .CK(clk), .Q(
        \xmem_inst/mem[3][0] ) );
  DFF_X1 \xmem_inst/mem_reg[3][1]  ( .D(n1265), .CK(clk), .Q(
        \xmem_inst/mem[3][1] ) );
  DFF_X1 \xmem_inst/mem_reg[3][2]  ( .D(n1264), .CK(clk), .Q(
        \xmem_inst/mem[3][2] ) );
  DFF_X1 \xmem_inst/mem_reg[3][3]  ( .D(n1263), .CK(clk), .Q(
        \xmem_inst/mem[3][3] ) );
  DFF_X1 \xmem_inst/mem_reg[3][4]  ( .D(n1262), .CK(clk), .Q(
        \xmem_inst/mem[3][4] ) );
  DFF_X1 \xmem_inst/mem_reg[3][5]  ( .D(n1261), .CK(clk), .Q(
        \xmem_inst/mem[3][5] ) );
  DFF_X1 \xmem_inst/mem_reg[3][6]  ( .D(n1260), .CK(clk), .Q(
        \xmem_inst/mem[3][6] ) );
  DFF_X1 \xmem_inst/mem_reg[3][7]  ( .D(n1259), .CK(clk), .Q(
        \xmem_inst/mem[3][7] ) );
  DFF_X1 \xmem_inst/mem_reg[3][8]  ( .D(n1258), .CK(clk), .Q(
        \xmem_inst/mem[3][8] ) );
  DFF_X1 \xmem_inst/mem_reg[3][9]  ( .D(n1257), .CK(clk), .Q(
        \xmem_inst/mem[3][9] ) );
  DFF_X1 \xmem_inst/mem_reg[3][10]  ( .D(n1256), .CK(clk), .Q(
        \xmem_inst/mem[3][10] ) );
  DFF_X1 \xmem_inst/mem_reg[3][11]  ( .D(n1255), .CK(clk), .Q(
        \xmem_inst/mem[3][11] ) );
  DFF_X1 \xmem_inst/mem_reg[3][12]  ( .D(n1254), .CK(clk), .Q(
        \xmem_inst/mem[3][12] ) );
  DFF_X1 \xmem_inst/mem_reg[3][13]  ( .D(n1253), .CK(clk), .Q(
        \xmem_inst/mem[3][13] ) );
  DFF_X1 \xmem_inst/mem_reg[3][14]  ( .D(n1252), .CK(clk), .Q(
        \xmem_inst/mem[3][14] ) );
  DFF_X1 \xmem_inst/mem_reg[3][15]  ( .D(n1251), .CK(clk), .Q(
        \xmem_inst/mem[3][15] ) );
  DFF_X1 \xmem_inst/mem_reg[3][16]  ( .D(n1250), .CK(clk), .Q(
        \xmem_inst/mem[3][16] ) );
  DFF_X1 \xmem_inst/mem_reg[3][17]  ( .D(n1249), .CK(clk), .Q(
        \xmem_inst/mem[3][17] ) );
  DFF_X1 \xmem_inst/mem_reg[3][18]  ( .D(n1248), .CK(clk), .Q(
        \xmem_inst/mem[3][18] ) );
  DFF_X1 \xmem_inst/mem_reg[3][19]  ( .D(n1247), .CK(clk), .Q(
        \xmem_inst/mem[3][19] ) );
  DFF_X1 \xmem_inst/mem_reg[4][0]  ( .D(n1246), .CK(clk), .Q(
        \xmem_inst/mem[4][0] ) );
  DFF_X1 \xmem_inst/mem_reg[4][1]  ( .D(n1245), .CK(clk), .Q(
        \xmem_inst/mem[4][1] ) );
  DFF_X1 \xmem_inst/mem_reg[4][2]  ( .D(n1244), .CK(clk), .Q(
        \xmem_inst/mem[4][2] ) );
  DFF_X1 \xmem_inst/mem_reg[4][3]  ( .D(n1243), .CK(clk), .Q(
        \xmem_inst/mem[4][3] ) );
  DFF_X1 \xmem_inst/mem_reg[4][4]  ( .D(n1242), .CK(clk), .Q(
        \xmem_inst/mem[4][4] ) );
  DFF_X1 \xmem_inst/mem_reg[4][5]  ( .D(n1241), .CK(clk), .Q(
        \xmem_inst/mem[4][5] ) );
  DFF_X1 \xmem_inst/mem_reg[4][6]  ( .D(n1240), .CK(clk), .Q(
        \xmem_inst/mem[4][6] ) );
  DFF_X1 \xmem_inst/mem_reg[4][7]  ( .D(n1239), .CK(clk), .Q(
        \xmem_inst/mem[4][7] ) );
  DFF_X1 \xmem_inst/mem_reg[4][8]  ( .D(n1238), .CK(clk), .Q(
        \xmem_inst/mem[4][8] ) );
  DFF_X1 \xmem_inst/mem_reg[4][9]  ( .D(n1237), .CK(clk), .Q(
        \xmem_inst/mem[4][9] ) );
  DFF_X1 \xmem_inst/mem_reg[4][10]  ( .D(n1236), .CK(clk), .Q(
        \xmem_inst/mem[4][10] ) );
  DFF_X1 \xmem_inst/mem_reg[4][11]  ( .D(n1235), .CK(clk), .Q(
        \xmem_inst/mem[4][11] ) );
  DFF_X1 \xmem_inst/mem_reg[4][12]  ( .D(n1234), .CK(clk), .Q(
        \xmem_inst/mem[4][12] ) );
  DFF_X1 \xmem_inst/mem_reg[4][13]  ( .D(n1233), .CK(clk), .Q(
        \xmem_inst/mem[4][13] ) );
  DFF_X1 \xmem_inst/mem_reg[4][14]  ( .D(n1232), .CK(clk), .Q(
        \xmem_inst/mem[4][14] ) );
  DFF_X1 \xmem_inst/mem_reg[4][15]  ( .D(n1231), .CK(clk), .Q(
        \xmem_inst/mem[4][15] ) );
  DFF_X1 \xmem_inst/mem_reg[4][16]  ( .D(n1230), .CK(clk), .Q(
        \xmem_inst/mem[4][16] ) );
  DFF_X1 \xmem_inst/mem_reg[4][17]  ( .D(n1229), .CK(clk), .Q(
        \xmem_inst/mem[4][17] ) );
  DFF_X1 \xmem_inst/mem_reg[4][18]  ( .D(n1228), .CK(clk), .Q(
        \xmem_inst/mem[4][18] ) );
  DFF_X1 \xmem_inst/mem_reg[4][19]  ( .D(n1227), .CK(clk), .Q(
        \xmem_inst/mem[4][19] ) );
  DFF_X1 \xmem_inst/mem_reg[5][0]  ( .D(n1226), .CK(clk), .Q(
        \xmem_inst/mem[5][0] ) );
  DFF_X1 \xmem_inst/mem_reg[5][1]  ( .D(n1225), .CK(clk), .Q(
        \xmem_inst/mem[5][1] ) );
  DFF_X1 \xmem_inst/mem_reg[5][2]  ( .D(n1224), .CK(clk), .Q(
        \xmem_inst/mem[5][2] ) );
  DFF_X1 \xmem_inst/mem_reg[5][3]  ( .D(n1223), .CK(clk), .Q(
        \xmem_inst/mem[5][3] ) );
  DFF_X1 \xmem_inst/mem_reg[5][4]  ( .D(n1222), .CK(clk), .Q(
        \xmem_inst/mem[5][4] ) );
  DFF_X1 \xmem_inst/mem_reg[5][5]  ( .D(n1221), .CK(clk), .Q(
        \xmem_inst/mem[5][5] ) );
  DFF_X1 \xmem_inst/mem_reg[5][6]  ( .D(n1220), .CK(clk), .Q(
        \xmem_inst/mem[5][6] ) );
  DFF_X1 \xmem_inst/mem_reg[5][7]  ( .D(n1219), .CK(clk), .Q(
        \xmem_inst/mem[5][7] ) );
  DFF_X1 \xmem_inst/mem_reg[5][8]  ( .D(n1218), .CK(clk), .Q(
        \xmem_inst/mem[5][8] ) );
  DFF_X1 \xmem_inst/mem_reg[5][9]  ( .D(n1217), .CK(clk), .Q(
        \xmem_inst/mem[5][9] ) );
  DFF_X1 \xmem_inst/mem_reg[5][10]  ( .D(n1216), .CK(clk), .Q(
        \xmem_inst/mem[5][10] ) );
  DFF_X1 \xmem_inst/mem_reg[5][11]  ( .D(n1215), .CK(clk), .Q(
        \xmem_inst/mem[5][11] ) );
  DFF_X1 \xmem_inst/mem_reg[5][12]  ( .D(n1214), .CK(clk), .Q(
        \xmem_inst/mem[5][12] ) );
  DFF_X1 \xmem_inst/mem_reg[5][13]  ( .D(n1213), .CK(clk), .Q(
        \xmem_inst/mem[5][13] ) );
  DFF_X1 \xmem_inst/mem_reg[5][14]  ( .D(n1212), .CK(clk), .Q(
        \xmem_inst/mem[5][14] ) );
  DFF_X1 \xmem_inst/mem_reg[5][15]  ( .D(n1211), .CK(clk), .Q(
        \xmem_inst/mem[5][15] ) );
  DFF_X1 \xmem_inst/mem_reg[5][16]  ( .D(n1210), .CK(clk), .Q(
        \xmem_inst/mem[5][16] ) );
  DFF_X1 \xmem_inst/mem_reg[5][17]  ( .D(n1209), .CK(clk), .Q(
        \xmem_inst/mem[5][17] ) );
  DFF_X1 \xmem_inst/mem_reg[5][18]  ( .D(n1208), .CK(clk), .Q(
        \xmem_inst/mem[5][18] ) );
  DFF_X1 \xmem_inst/mem_reg[5][19]  ( .D(n1207), .CK(clk), .Q(
        \xmem_inst/mem[5][19] ) );
  DFF_X1 \xmem_inst/mem_reg[6][0]  ( .D(n1206), .CK(clk), .Q(
        \xmem_inst/mem[6][0] ) );
  DFF_X1 \xmem_inst/mem_reg[6][1]  ( .D(n1205), .CK(clk), .Q(
        \xmem_inst/mem[6][1] ) );
  DFF_X1 \xmem_inst/mem_reg[6][2]  ( .D(n1204), .CK(clk), .Q(
        \xmem_inst/mem[6][2] ) );
  DFF_X1 \xmem_inst/mem_reg[6][3]  ( .D(n1203), .CK(clk), .Q(
        \xmem_inst/mem[6][3] ) );
  DFF_X1 \xmem_inst/mem_reg[6][4]  ( .D(n1202), .CK(clk), .Q(
        \xmem_inst/mem[6][4] ) );
  DFF_X1 \xmem_inst/mem_reg[6][5]  ( .D(n1201), .CK(clk), .Q(
        \xmem_inst/mem[6][5] ) );
  DFF_X1 \xmem_inst/mem_reg[6][6]  ( .D(n1200), .CK(clk), .Q(
        \xmem_inst/mem[6][6] ) );
  DFF_X1 \xmem_inst/mem_reg[6][7]  ( .D(n1199), .CK(clk), .Q(
        \xmem_inst/mem[6][7] ) );
  DFF_X1 \xmem_inst/mem_reg[6][8]  ( .D(n1198), .CK(clk), .Q(
        \xmem_inst/mem[6][8] ) );
  DFF_X1 \xmem_inst/mem_reg[6][9]  ( .D(n1197), .CK(clk), .Q(
        \xmem_inst/mem[6][9] ) );
  DFF_X1 \xmem_inst/mem_reg[6][10]  ( .D(n1196), .CK(clk), .Q(
        \xmem_inst/mem[6][10] ) );
  DFF_X1 \xmem_inst/mem_reg[6][11]  ( .D(n1195), .CK(clk), .Q(
        \xmem_inst/mem[6][11] ) );
  DFF_X1 \xmem_inst/mem_reg[6][12]  ( .D(n1194), .CK(clk), .Q(
        \xmem_inst/mem[6][12] ) );
  DFF_X1 \xmem_inst/mem_reg[6][13]  ( .D(n1193), .CK(clk), .Q(
        \xmem_inst/mem[6][13] ) );
  DFF_X1 \xmem_inst/mem_reg[6][14]  ( .D(n1192), .CK(clk), .Q(
        \xmem_inst/mem[6][14] ) );
  DFF_X1 \xmem_inst/mem_reg[6][15]  ( .D(n1191), .CK(clk), .Q(
        \xmem_inst/mem[6][15] ) );
  DFF_X1 \xmem_inst/mem_reg[6][16]  ( .D(n1190), .CK(clk), .Q(
        \xmem_inst/mem[6][16] ) );
  DFF_X1 \xmem_inst/mem_reg[6][17]  ( .D(n1189), .CK(clk), .Q(
        \xmem_inst/mem[6][17] ) );
  DFF_X1 \xmem_inst/mem_reg[6][18]  ( .D(n1188), .CK(clk), .Q(
        \xmem_inst/mem[6][18] ) );
  DFF_X1 \xmem_inst/mem_reg[6][19]  ( .D(n1187), .CK(clk), .Q(
        \xmem_inst/mem[6][19] ) );
  DFF_X1 \xmem_inst/mem_reg[7][0]  ( .D(n1186), .CK(clk), .Q(
        \xmem_inst/mem[7][0] ) );
  DFF_X1 \xmem_inst/mem_reg[7][1]  ( .D(n1185), .CK(clk), .Q(
        \xmem_inst/mem[7][1] ) );
  DFF_X1 \xmem_inst/mem_reg[7][2]  ( .D(n1184), .CK(clk), .Q(
        \xmem_inst/mem[7][2] ) );
  DFF_X1 \xmem_inst/mem_reg[7][3]  ( .D(n1183), .CK(clk), .Q(
        \xmem_inst/mem[7][3] ) );
  DFF_X1 \xmem_inst/mem_reg[7][4]  ( .D(n1182), .CK(clk), .Q(
        \xmem_inst/mem[7][4] ) );
  DFF_X1 \xmem_inst/mem_reg[7][5]  ( .D(n1181), .CK(clk), .Q(
        \xmem_inst/mem[7][5] ) );
  DFF_X1 \xmem_inst/mem_reg[7][6]  ( .D(n1180), .CK(clk), .Q(
        \xmem_inst/mem[7][6] ) );
  DFF_X1 \xmem_inst/mem_reg[7][7]  ( .D(n1179), .CK(clk), .Q(
        \xmem_inst/mem[7][7] ) );
  DFF_X1 \xmem_inst/mem_reg[7][8]  ( .D(n1178), .CK(clk), .Q(
        \xmem_inst/mem[7][8] ) );
  DFF_X1 \xmem_inst/mem_reg[7][9]  ( .D(n1177), .CK(clk), .Q(
        \xmem_inst/mem[7][9] ) );
  DFF_X1 \xmem_inst/mem_reg[7][10]  ( .D(n1176), .CK(clk), .Q(
        \xmem_inst/mem[7][10] ) );
  DFF_X1 \xmem_inst/mem_reg[7][11]  ( .D(n1175), .CK(clk), .Q(
        \xmem_inst/mem[7][11] ) );
  DFF_X1 \xmem_inst/mem_reg[7][12]  ( .D(n1174), .CK(clk), .Q(
        \xmem_inst/mem[7][12] ) );
  DFF_X1 \xmem_inst/mem_reg[7][13]  ( .D(n1173), .CK(clk), .Q(
        \xmem_inst/mem[7][13] ) );
  DFF_X1 \xmem_inst/mem_reg[7][14]  ( .D(n1172), .CK(clk), .Q(
        \xmem_inst/mem[7][14] ) );
  DFF_X1 \xmem_inst/mem_reg[7][15]  ( .D(n1171), .CK(clk), .Q(
        \xmem_inst/mem[7][15] ) );
  DFF_X1 \xmem_inst/mem_reg[7][16]  ( .D(n1170), .CK(clk), .Q(
        \xmem_inst/mem[7][16] ) );
  DFF_X1 \xmem_inst/mem_reg[7][17]  ( .D(n1169), .CK(clk), .Q(
        \xmem_inst/mem[7][17] ) );
  DFF_X1 \xmem_inst/mem_reg[7][18]  ( .D(n1168), .CK(clk), .Q(
        \xmem_inst/mem[7][18] ) );
  DFF_X1 \xmem_inst/mem_reg[7][19]  ( .D(n1167), .CK(clk), .Q(
        \xmem_inst/mem[7][19] ) );
  DFF_X1 \xmem_inst/mem_reg[16][0]  ( .D(n1006), .CK(clk), .Q(
        \xmem_inst/mem[16][0] ) );
  DFF_X1 \xmem_inst/mem_reg[16][1]  ( .D(n1005), .CK(clk), .Q(
        \xmem_inst/mem[16][1] ) );
  DFF_X1 \xmem_inst/mem_reg[16][2]  ( .D(n1004), .CK(clk), .Q(
        \xmem_inst/mem[16][2] ) );
  DFF_X1 \xmem_inst/mem_reg[16][3]  ( .D(n1003), .CK(clk), .Q(
        \xmem_inst/mem[16][3] ) );
  DFF_X1 \xmem_inst/mem_reg[16][4]  ( .D(n1002), .CK(clk), .Q(
        \xmem_inst/mem[16][4] ) );
  DFF_X1 \xmem_inst/mem_reg[16][5]  ( .D(n1001), .CK(clk), .Q(
        \xmem_inst/mem[16][5] ) );
  DFF_X1 \xmem_inst/mem_reg[16][6]  ( .D(n1000), .CK(clk), .Q(
        \xmem_inst/mem[16][6] ) );
  DFF_X1 \xmem_inst/mem_reg[16][7]  ( .D(n999), .CK(clk), .Q(
        \xmem_inst/mem[16][7] ) );
  DFF_X1 \xmem_inst/mem_reg[16][8]  ( .D(n998), .CK(clk), .Q(
        \xmem_inst/mem[16][8] ) );
  DFF_X1 \xmem_inst/mem_reg[16][9]  ( .D(n997), .CK(clk), .Q(
        \xmem_inst/mem[16][9] ) );
  DFF_X1 \xmem_inst/mem_reg[16][10]  ( .D(n996), .CK(clk), .Q(
        \xmem_inst/mem[16][10] ) );
  DFF_X1 \xmem_inst/mem_reg[16][11]  ( .D(n995), .CK(clk), .Q(
        \xmem_inst/mem[16][11] ) );
  DFF_X1 \xmem_inst/mem_reg[16][12]  ( .D(n994), .CK(clk), .Q(
        \xmem_inst/mem[16][12] ) );
  DFF_X1 \xmem_inst/mem_reg[16][13]  ( .D(n993), .CK(clk), .Q(
        \xmem_inst/mem[16][13] ) );
  DFF_X1 \xmem_inst/mem_reg[16][14]  ( .D(n992), .CK(clk), .Q(
        \xmem_inst/mem[16][14] ) );
  DFF_X1 \xmem_inst/mem_reg[16][15]  ( .D(n991), .CK(clk), .Q(
        \xmem_inst/mem[16][15] ) );
  DFF_X1 \xmem_inst/mem_reg[16][16]  ( .D(n990), .CK(clk), .Q(
        \xmem_inst/mem[16][16] ) );
  DFF_X1 \xmem_inst/mem_reg[16][17]  ( .D(n989), .CK(clk), .Q(
        \xmem_inst/mem[16][17] ) );
  DFF_X1 \xmem_inst/mem_reg[16][18]  ( .D(n988), .CK(clk), .Q(
        \xmem_inst/mem[16][18] ) );
  DFF_X1 \xmem_inst/mem_reg[16][19]  ( .D(n987), .CK(clk), .Q(
        \xmem_inst/mem[16][19] ) );
  DFF_X1 \xmem_inst/mem_reg[17][0]  ( .D(n986), .CK(clk), .Q(
        \xmem_inst/mem[17][0] ) );
  DFF_X1 \xmem_inst/mem_reg[17][1]  ( .D(n985), .CK(clk), .Q(
        \xmem_inst/mem[17][1] ) );
  DFF_X1 \xmem_inst/mem_reg[17][2]  ( .D(n984), .CK(clk), .Q(
        \xmem_inst/mem[17][2] ) );
  DFF_X1 \xmem_inst/mem_reg[17][3]  ( .D(n983), .CK(clk), .Q(
        \xmem_inst/mem[17][3] ) );
  DFF_X1 \xmem_inst/mem_reg[17][4]  ( .D(n982), .CK(clk), .Q(
        \xmem_inst/mem[17][4] ) );
  DFF_X1 \xmem_inst/mem_reg[17][5]  ( .D(n981), .CK(clk), .Q(
        \xmem_inst/mem[17][5] ) );
  DFF_X1 \xmem_inst/mem_reg[17][6]  ( .D(n980), .CK(clk), .Q(
        \xmem_inst/mem[17][6] ) );
  DFF_X1 \xmem_inst/mem_reg[17][7]  ( .D(n979), .CK(clk), .Q(
        \xmem_inst/mem[17][7] ) );
  DFF_X1 \xmem_inst/mem_reg[17][8]  ( .D(n978), .CK(clk), .Q(
        \xmem_inst/mem[17][8] ) );
  DFF_X1 \xmem_inst/mem_reg[17][9]  ( .D(n977), .CK(clk), .Q(
        \xmem_inst/mem[17][9] ) );
  DFF_X1 \xmem_inst/mem_reg[17][10]  ( .D(n976), .CK(clk), .Q(
        \xmem_inst/mem[17][10] ) );
  DFF_X1 \xmem_inst/mem_reg[17][11]  ( .D(n975), .CK(clk), .Q(
        \xmem_inst/mem[17][11] ) );
  DFF_X1 \xmem_inst/mem_reg[17][12]  ( .D(n974), .CK(clk), .Q(
        \xmem_inst/mem[17][12] ) );
  DFF_X1 \xmem_inst/mem_reg[17][13]  ( .D(n973), .CK(clk), .Q(
        \xmem_inst/mem[17][13] ) );
  DFF_X1 \xmem_inst/mem_reg[17][14]  ( .D(n972), .CK(clk), .Q(
        \xmem_inst/mem[17][14] ) );
  DFF_X1 \xmem_inst/mem_reg[17][15]  ( .D(n971), .CK(clk), .Q(
        \xmem_inst/mem[17][15] ) );
  DFF_X1 \xmem_inst/mem_reg[17][16]  ( .D(n970), .CK(clk), .Q(
        \xmem_inst/mem[17][16] ) );
  DFF_X1 \xmem_inst/mem_reg[17][17]  ( .D(n969), .CK(clk), .Q(
        \xmem_inst/mem[17][17] ) );
  DFF_X1 \xmem_inst/mem_reg[17][18]  ( .D(n968), .CK(clk), .Q(
        \xmem_inst/mem[17][18] ) );
  DFF_X1 \xmem_inst/mem_reg[17][19]  ( .D(n967), .CK(clk), .Q(
        \xmem_inst/mem[17][19] ) );
  DFF_X1 \xmem_inst/mem_reg[18][0]  ( .D(n966), .CK(clk), .Q(
        \xmem_inst/mem[18][0] ) );
  DFF_X1 \xmem_inst/mem_reg[18][1]  ( .D(n965), .CK(clk), .Q(
        \xmem_inst/mem[18][1] ) );
  DFF_X1 \xmem_inst/mem_reg[18][2]  ( .D(n964), .CK(clk), .Q(
        \xmem_inst/mem[18][2] ) );
  DFF_X1 \xmem_inst/mem_reg[18][3]  ( .D(n963), .CK(clk), .Q(
        \xmem_inst/mem[18][3] ) );
  DFF_X1 \xmem_inst/mem_reg[18][4]  ( .D(n962), .CK(clk), .Q(
        \xmem_inst/mem[18][4] ) );
  DFF_X1 \xmem_inst/mem_reg[18][5]  ( .D(n961), .CK(clk), .Q(
        \xmem_inst/mem[18][5] ) );
  DFF_X1 \xmem_inst/mem_reg[18][6]  ( .D(n960), .CK(clk), .Q(
        \xmem_inst/mem[18][6] ) );
  DFF_X1 \xmem_inst/mem_reg[18][7]  ( .D(n959), .CK(clk), .Q(
        \xmem_inst/mem[18][7] ) );
  DFF_X1 \xmem_inst/mem_reg[18][8]  ( .D(n958), .CK(clk), .Q(
        \xmem_inst/mem[18][8] ) );
  DFF_X1 \xmem_inst/mem_reg[18][9]  ( .D(n957), .CK(clk), .Q(
        \xmem_inst/mem[18][9] ) );
  DFF_X1 \xmem_inst/mem_reg[18][10]  ( .D(n956), .CK(clk), .Q(
        \xmem_inst/mem[18][10] ) );
  DFF_X1 \xmem_inst/mem_reg[18][11]  ( .D(n955), .CK(clk), .Q(
        \xmem_inst/mem[18][11] ) );
  DFF_X1 \xmem_inst/mem_reg[18][12]  ( .D(n954), .CK(clk), .Q(
        \xmem_inst/mem[18][12] ) );
  DFF_X1 \xmem_inst/mem_reg[18][13]  ( .D(n953), .CK(clk), .Q(
        \xmem_inst/mem[18][13] ) );
  DFF_X1 \xmem_inst/mem_reg[18][14]  ( .D(n952), .CK(clk), .Q(
        \xmem_inst/mem[18][14] ) );
  DFF_X1 \xmem_inst/mem_reg[18][15]  ( .D(n951), .CK(clk), .Q(
        \xmem_inst/mem[18][15] ) );
  DFF_X1 \xmem_inst/mem_reg[18][16]  ( .D(n950), .CK(clk), .Q(
        \xmem_inst/mem[18][16] ) );
  DFF_X1 \xmem_inst/mem_reg[18][17]  ( .D(n949), .CK(clk), .Q(
        \xmem_inst/mem[18][17] ) );
  DFF_X1 \xmem_inst/mem_reg[18][18]  ( .D(n948), .CK(clk), .Q(
        \xmem_inst/mem[18][18] ) );
  DFF_X1 \xmem_inst/mem_reg[18][19]  ( .D(n947), .CK(clk), .Q(
        \xmem_inst/mem[18][19] ) );
  DFF_X1 \fmem_addr_reg[0]  ( .D(n926), .CK(clk), .Q(fmem_addr[0]), .QN(n3331)
         );
  DFF_X1 \fmem_addr_reg[2]  ( .D(n924), .CK(clk), .Q(fmem_addr[2]), .QN(n3332)
         );
  DFF_X1 \xmem_inst/mem_reg[19][0]  ( .D(n946), .CK(clk), .Q(
        \xmem_inst/mem[19][0] ) );
  DFF_X1 \xmem_inst/mem_reg[19][1]  ( .D(n945), .CK(clk), .Q(
        \xmem_inst/mem[19][1] ) );
  DFF_X1 \xmem_inst/mem_reg[19][2]  ( .D(n944), .CK(clk), .Q(
        \xmem_inst/mem[19][2] ) );
  DFF_X1 \xmem_inst/data_out_reg[2]  ( .D(\xmem_inst/N107 ), .CK(clk), .Q(
        xmem_data[2]), .QN(n1345) );
  DFF_X1 \xmem_inst/mem_reg[19][3]  ( .D(n943), .CK(clk), .Q(
        \xmem_inst/mem[19][3] ) );
  DFF_X1 \xmem_inst/mem_reg[19][4]  ( .D(n942), .CK(clk), .Q(
        \xmem_inst/mem[19][4] ) );
  DFF_X1 \xmem_inst/data_out_reg[4]  ( .D(\xmem_inst/N105 ), .CK(clk), .Q(
        xmem_data[4]) );
  DFF_X1 \xmem_inst/mem_reg[19][5]  ( .D(n941), .CK(clk), .Q(
        \xmem_inst/mem[19][5] ) );
  DFF_X1 \xmem_inst/mem_reg[19][6]  ( .D(n940), .CK(clk), .Q(
        \xmem_inst/mem[19][6] ) );
  DFF_X1 \xmem_inst/data_out_reg[6]  ( .D(\xmem_inst/N103 ), .CK(clk), .Q(
        xmem_data[6]), .QN(n3317) );
  DFF_X1 \xmem_inst/mem_reg[19][7]  ( .D(n939), .CK(clk), .Q(
        \xmem_inst/mem[19][7] ) );
  DFF_X1 \xmem_inst/mem_reg[19][8]  ( .D(n938), .CK(clk), .Q(
        \xmem_inst/mem[19][8] ) );
  DFF_X1 \xmem_inst/data_out_reg[8]  ( .D(\xmem_inst/N101 ), .CK(clk), .Q(
        xmem_data[8]) );
  DFF_X1 \xmem_inst/mem_reg[19][9]  ( .D(n937), .CK(clk), .Q(
        \xmem_inst/mem[19][9] ) );
  DFF_X1 \xmem_inst/mem_reg[19][10]  ( .D(n936), .CK(clk), .Q(
        \xmem_inst/mem[19][10] ) );
  DFF_X1 \xmem_inst/data_out_reg[10]  ( .D(\xmem_inst/N99 ), .CK(clk), .Q(
        xmem_data[10]), .QN(n3323) );
  DFF_X1 \xmem_inst/mem_reg[19][11]  ( .D(n935), .CK(clk), .Q(
        \xmem_inst/mem[19][11] ) );
  DFF_X1 \xmem_inst/mem_reg[19][12]  ( .D(n934), .CK(clk), .Q(
        \xmem_inst/mem[19][12] ) );
  DFF_X1 \xmem_inst/data_out_reg[12]  ( .D(\xmem_inst/N97 ), .CK(clk), .Q(
        xmem_data[12]), .QN(n3319) );
  DFF_X1 \xmem_inst/mem_reg[19][13]  ( .D(n933), .CK(clk), .Q(
        \xmem_inst/mem[19][13] ) );
  DFF_X1 \xmem_inst/mem_reg[19][14]  ( .D(n932), .CK(clk), .Q(
        \xmem_inst/mem[19][14] ) );
  DFF_X1 \xmem_inst/data_out_reg[14]  ( .D(\xmem_inst/N95 ), .CK(clk), .Q(
        xmem_data[14]), .QN(n3316) );
  DFF_X1 \xmem_inst/mem_reg[19][15]  ( .D(n931), .CK(clk), .Q(
        \xmem_inst/mem[19][15] ) );
  DFF_X1 \xmem_inst/mem_reg[19][16]  ( .D(n930), .CK(clk), .Q(
        \xmem_inst/mem[19][16] ) );
  DFF_X1 \xmem_inst/data_out_reg[16]  ( .D(\xmem_inst/N93 ), .CK(clk), .Q(
        xmem_data[16]), .QN(n3315) );
  DFF_X1 \xmem_inst/mem_reg[19][17]  ( .D(n929), .CK(clk), .Q(
        \xmem_inst/mem[19][17] ) );
  DFF_X1 \xmem_inst/mem_reg[19][18]  ( .D(n928), .CK(clk), .Q(
        \xmem_inst/mem[19][18] ) );
  DFF_X1 \xmem_inst/mem_reg[19][19]  ( .D(n927), .CK(clk), .Q(
        \xmem_inst/mem[19][19] ) );
  DFF_X1 \ctrl_conv_output_inst/conv_start_accum_reg  ( .D(
        \ctrl_conv_output_inst/N74 ), .CK(clk), .Q(
        \ctrl_conv_output_inst/conv_start_accum ), .QN(n3368) );
  DFF_X1 \fmem_inst/z_reg[5]  ( .D(n917), .CK(clk), .Q(fmem_data[5]) );
  DFF_X1 \fmem_inst/z_reg[1]  ( .D(n921), .CK(clk), .Q(fmem_data[1]) );
  DFF_X1 \fmem_inst/z_reg[2]  ( .D(n920), .CK(clk), .Q(fmem_data[2]), .QN(
        n1346) );
  DFF_X1 \fmem_inst/z_reg[3]  ( .D(n919), .CK(clk), .Q(fmem_data[3]), .QN(
        n1349) );
  DFF_X1 \fmem_inst/z_reg[6]  ( .D(n916), .CK(clk), .Q(fmem_data[6]), .QN(
        n1347) );
  DFF_X1 \fmem_inst/z_reg[7]  ( .D(n915), .CK(clk), .Q(fmem_data[7]), .QN(
        n1350) );
  DFF_X1 \fmem_inst/z_reg[9]  ( .D(n913), .CK(clk), .Q(fmem_data[9]), .QN(
        n1348) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[0]  ( .D(n890), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [0]), .QN(n3348) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[1]  ( .D(n889), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [1]), .QN(n3349) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[2]  ( .D(n888), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [2]), .QN(n3350) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[3]  ( .D(n887), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [3]), .QN(n3351) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[4]  ( .D(n886), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [4]), .QN(n3352) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[5]  ( .D(n885), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [5]), .QN(n3353) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[6]  ( .D(n884), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [6]), .QN(n3354) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[7]  ( .D(n883), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [7]), .QN(n3355) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[8]  ( .D(n882), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [8]), .QN(n3356) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[9]  ( .D(n881), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [9]), .QN(n3357) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[10]  ( .D(n880), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [10]), .QN(n3358) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[11]  ( .D(n879), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [11]), .QN(n3364) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[12]  ( .D(n878), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [12]), .QN(n3359) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[13]  ( .D(n877), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [13]), .QN(n3360) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[14]  ( .D(n876), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [14]), .QN(n3361) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[15]  ( .D(n875), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [15]), .QN(n3362) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[16]  ( .D(n874), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [16]), .QN(n3363) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[17]  ( .D(n873), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [17]), .QN(n3365) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[18]  ( .D(n872), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [18]), .QN(n3366) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[19]  ( .D(n871), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [19]), .QN(n3369) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[0]  ( .D(n910), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [0]), .QN(n3378) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[1]  ( .D(n909), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [1]), .QN(n3379) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[3]  ( .D(n907), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [3]), .QN(n3370) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[4]  ( .D(n906), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [4]), .QN(n3381) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[5]  ( .D(n905), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [5]), .QN(n3371) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[6]  ( .D(n904), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [6]), .QN(n3382) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[7]  ( .D(n903), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [7]), .QN(n3372) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[8]  ( .D(n902), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [8]), .QN(n3383) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[9]  ( .D(n901), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [9]), .QN(n3373) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[10]  ( .D(n900), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [10]), .QN(n3384) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[11]  ( .D(n899), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [11]), .QN(n3374) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[12]  ( .D(n898), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [12]), .QN(n3385) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[14]  ( .D(n896), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [14]), .QN(n3386) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[15]  ( .D(n895), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [15]), .QN(n3376) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[17]  ( .D(n893), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [17]), .QN(n3377) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[19]  ( .D(n891), .CK(clk), .QN(n3325)
         );
  DFF_X1 \xmem_inst/data_out_reg[11]  ( .D(\xmem_inst/N98 ), .CK(clk), .Q(
        n3320), .QN(n3391) );
  DFF_X1 \fmem_addr_reg[1]  ( .D(n925), .CK(clk), .Q(fmem_addr[1]), .QN(n3347)
         );
  DFF_X1 \xmem_inst/data_out_reg[9]  ( .D(\xmem_inst/N100 ), .CK(clk), .Q(
        xmem_data[9]), .QN(n3322) );
  DFF_X1 \xmem_inst/data_out_reg[3]  ( .D(\xmem_inst/N106 ), .CK(clk), .Q(
        xmem_data[3]), .QN(n1352) );
  DFF_X1 \xmem_inst/data_out_reg[7]  ( .D(n1382), .CK(clk), .Q(n3329), .QN(
        xmem_data[7]) );
  DFF_X1 \xmem_inst/data_out_reg[5]  ( .D(n1381), .CK(clk), .Q(n3321), .QN(
        xmem_data[5]) );
  DFF_X1 \xmem_inst/data_out_reg[13]  ( .D(n1380), .CK(clk), .Q(n3327), .QN(
        \DP_OP_485J1_122_4413/n1657 ) );
  DFF_X1 \xmem_inst/data_out_reg[17]  ( .D(n1379), .CK(clk), .Q(n3318), .QN(
        \DP_OP_485J1_122_4413/n1655 ) );
  DFF_X1 \xmem_inst/data_out_reg[19]  ( .D(n1378), .CK(clk), .Q(n3326), .QN(
        xmem_data[19]) );
  DFF_X2 \fmem_inst/z_reg[19]  ( .D(n912), .CK(clk), .Q(fmem_data[19]) );
  SDFF_X1 \xmem_inst/data_out_reg[15]  ( .D(\xmem_inst/N94 ), .SI(1'b0), .SE(
        1'b0), .CK(clk), .Q(\DP_OP_485J1_122_4413/n1656 ), .QN(n1351) );
  DFF_X1 \xmem_inst/data_out_reg[18]  ( .D(\xmem_inst/N91 ), .CK(clk), .Q(
        xmem_data[18]), .QN(n3324) );
  DFF_X1 \xmem_inst/data_out_reg[0]  ( .D(\xmem_inst/N109 ), .CK(clk), .Q(
        xmem_data[0]), .QN(n3328) );
  DFF_X1 \fmem_inst/z_reg[4]  ( .D(n918), .CK(clk), .Q(fmem_data[4]), .QN(
        n3390) );
  DFF_X1 \fmem_inst/z_reg[8]  ( .D(n914), .CK(clk), .Q(fmem_data[8]), .QN(
        n3389) );
  DFFS_X1 \mac_unit_inst/x_mult_f_reg_reg[18]  ( .D(n892), .CK(clk), .SN(1'b1), 
        .Q(\mac_unit_inst/x_mult_f_reg [18]), .QN(n3388) );
  DFFS_X1 \mac_unit_inst/x_mult_f_reg_reg[16]  ( .D(n894), .CK(clk), .SN(1'b1), 
        .Q(\mac_unit_inst/x_mult_f_reg [16]), .QN(n3387) );
  DFFS_X1 \mac_unit_inst/x_mult_f_reg_reg[13]  ( .D(n897), .CK(clk), .SN(1'b1), 
        .Q(\mac_unit_inst/x_mult_f_reg [13]), .QN(n3375) );
  DFFS_X1 \mac_unit_inst/x_mult_f_reg_reg[2]  ( .D(n908), .CK(clk), .SN(1'b1), 
        .Q(\mac_unit_inst/x_mult_f_reg [2]), .QN(n3380) );
  SDFF_X2 \fmem_inst/z_reg[0]  ( .D(n922), .SI(1'b0), .SE(1'b0), .CK(clk), .Q(
        \DP_OP_485J1_122_4413/n1204 ), .QN(n3346) );
  DFF_X1 \xmem_inst/data_out_reg[1]  ( .D(n1384), .CK(clk), .Q(n3330), .QN(
        xmem_data[1]) );
  XOR2_X1 U1385 ( .A(n3330), .B(xmem_data[2]), .Z(n1882) );
  BUF_X1 U1386 ( .A(n1702), .Z(n1831) );
  INV_X1 U1387 ( .A(n2175), .ZN(n1340) );
  NAND2_X1 U1388 ( .A1(n2652), .A2(n2651), .ZN(n2783) );
  OR2_X1 U1389 ( .A1(n1823), .A2(n1822), .ZN(n2186) );
  INV_X1 U1390 ( .A(n2974), .ZN(n2975) );
  INV_X1 U1391 ( .A(n3090), .ZN(n3110) );
  INV_X1 U1392 ( .A(n3228), .ZN(n3227) );
  INV_X1 U1393 ( .A(n3204), .ZN(n3205) );
  INV_X1 U1394 ( .A(n3019), .ZN(n3020) );
  INV_X1 U1395 ( .A(n3067), .ZN(n3087) );
  INV_X1 U1396 ( .A(n3045), .ZN(n3065) );
  INV_X1 U1397 ( .A(n2996), .ZN(n2997) );
  INV_X1 U1398 ( .A(n3297), .ZN(n3296) );
  INV_X1 U1399 ( .A(n3251), .ZN(n3250) );
  INV_X1 U1400 ( .A(n2906), .ZN(n2905) );
  INV_X1 U1401 ( .A(n3180), .ZN(n3181) );
  INV_X1 U1402 ( .A(n3157), .ZN(n3158) );
  INV_X1 U1403 ( .A(n2861), .ZN(n2860) );
  INV_X1 U1404 ( .A(n3042), .ZN(n3043) );
  INV_X1 U1405 ( .A(n2883), .ZN(n2882) );
  INV_X1 U1406 ( .A(n3134), .ZN(n3135) );
  INV_X1 U1407 ( .A(n3275), .ZN(n3274) );
  INV_X1 U1408 ( .A(n2929), .ZN(n2928) );
  INV_X1 U1409 ( .A(n2952), .ZN(n2953) );
  NAND2_X1 U1410 ( .A1(n2908), .A2(n2415), .ZN(n2861) );
  NAND2_X1 U1411 ( .A1(n2908), .A2(n2885), .ZN(n2906) );
  NAND2_X1 U1412 ( .A1(n2908), .A2(n2442), .ZN(n2929) );
  NAND2_X1 U1413 ( .A1(n3254), .A2(n3207), .ZN(n3228) );
  NAND2_X1 U1414 ( .A1(n2908), .A2(n2457), .ZN(n2883) );
  NAND2_X1 U1415 ( .A1(n3254), .A2(n2447), .ZN(n3297) );
  BUF_X1 U1416 ( .A(n1750), .Z(n1911) );
  NAND2_X1 U1417 ( .A1(n3254), .A2(n3230), .ZN(n3251) );
  NAND2_X1 U1418 ( .A1(n3254), .A2(n3253), .ZN(n3275) );
  NOR2_X2 U1419 ( .A1(n3184), .A2(n2213), .ZN(n2203) );
  NOR2_X2 U1420 ( .A1(n3114), .A2(n2215), .ZN(n2216) );
  NOR2_X2 U1421 ( .A1(n2213), .A2(n3160), .ZN(n2214) );
  NOR2_X2 U1422 ( .A1(n3137), .A2(n2215), .ZN(n2212) );
  NOR2_X2 U1423 ( .A1(n2213), .A2(n3114), .ZN(n2200) );
  NOR2_X2 U1424 ( .A1(n3114), .A2(n2206), .ZN(n2207) );
  NOR2_X2 U1425 ( .A1(n3137), .A2(n2206), .ZN(n2201) );
  NOR2_X2 U1426 ( .A1(n3160), .A2(n2206), .ZN(n2205) );
  NOR2_X2 U1427 ( .A1(n2215), .A2(n3160), .ZN(n2202) );
  NOR2_X2 U1428 ( .A1(n3137), .A2(n2213), .ZN(n2204) );
  INV_X1 U1429 ( .A(n1389), .ZN(n1546) );
  INV_X1 U1430 ( .A(n1391), .ZN(n1629) );
  NAND2_X1 U1431 ( .A1(n1743), .A2(n2031), .ZN(n2034) );
  NAND2_X1 U1432 ( .A1(n1947), .A2(n1948), .ZN(n1954) );
  INV_X1 U1433 ( .A(n1996), .ZN(n1734) );
  INV_X1 U1434 ( .A(n1997), .ZN(n1735) );
  OAI21_X1 U1435 ( .B1(n1707), .B2(n1706), .A(n1705), .ZN(n1740) );
  NAND2_X1 U1436 ( .A1(n1714), .A2(n1713), .ZN(n1705) );
  NOR2_X1 U1437 ( .A1(n1714), .A2(n1713), .ZN(n1707) );
  INV_X1 U1438 ( .A(n1715), .ZN(n1706) );
  XNOR2_X1 U1439 ( .A(n1689), .B(n1688), .ZN(n1742) );
  XNOR2_X1 U1440 ( .A(n1687), .B(n1686), .ZN(n1688) );
  XNOR2_X1 U1441 ( .A(n1716), .B(n1715), .ZN(n1998) );
  XNOR2_X1 U1442 ( .A(n1475), .B(n1474), .ZN(n1477) );
  XNOR2_X1 U1443 ( .A(n1815), .B(n1814), .ZN(n1820) );
  XNOR2_X1 U1444 ( .A(n1813), .B(n1812), .ZN(n1814) );
  NAND2_X1 U1445 ( .A1(n1786), .A2(n1785), .ZN(n1810) );
  OAI21_X1 U1446 ( .B1(n1790), .B2(n1787), .A(n1788), .ZN(n1786) );
  NAND2_X1 U1447 ( .A1(n1790), .A2(n1787), .ZN(n1785) );
  CLKBUF_X1 U1448 ( .A(n2150), .Z(n2312) );
  OR2_X1 U1449 ( .A1(n3307), .A2(n2165), .ZN(n2800) );
  INV_X1 U1450 ( .A(n3326), .ZN(n1607) );
  INV_X1 U1451 ( .A(n1948), .ZN(n1950) );
  BUF_X2 U1452 ( .A(xmem_data[9]), .Z(n1837) );
  BUF_X1 U1453 ( .A(n1546), .Z(n1601) );
  NAND2_X1 U1454 ( .A1(n1453), .A2(n1452), .ZN(n1407) );
  INV_X1 U1455 ( .A(n1973), .ZN(n1969) );
  XNOR2_X1 U1456 ( .A(n1879), .B(n1878), .ZN(n1952) );
  OR2_X1 U1457 ( .A1(n1871), .A2(n1870), .ZN(n1872) );
  CLKBUF_X1 U1458 ( .A(n2096), .Z(n2091) );
  XNOR2_X1 U1459 ( .A(n1980), .B(n1961), .ZN(n1990) );
  NOR2_X1 U1460 ( .A1(n1523), .A2(n1522), .ZN(n1526) );
  NAND2_X1 U1461 ( .A1(n1523), .A2(n1522), .ZN(n1524) );
  NAND2_X1 U1462 ( .A1(n1479), .A2(n1478), .ZN(n1446) );
  NAND2_X1 U1463 ( .A1(n1687), .A2(n1686), .ZN(n1671) );
  XNOR2_X1 U1464 ( .A(n1862), .B(n1861), .ZN(n1842) );
  NAND2_X1 U1465 ( .A1(n1848), .A2(n1847), .ZN(n1931) );
  NAND2_X1 U1466 ( .A1(n1846), .A2(n1845), .ZN(n1847) );
  NAND2_X1 U1467 ( .A1(n1844), .A2(n1843), .ZN(n1848) );
  OR2_X1 U1468 ( .A1(n1846), .A2(n1845), .ZN(n1843) );
  BUF_X2 U1469 ( .A(n1626), .Z(n1909) );
  XNOR2_X1 U1470 ( .A(n3330), .B(xmem_data[2]), .ZN(n1799) );
  AND2_X1 U1471 ( .A1(n1617), .A2(n1616), .ZN(n2063) );
  XOR2_X1 U1472 ( .A(n2129), .B(n2128), .Z(n1616) );
  NAND2_X1 U1473 ( .A1(n1712), .A2(n1711), .ZN(n2153) );
  NAND2_X1 U1474 ( .A1(n1740), .A2(n1739), .ZN(n1711) );
  NAND2_X1 U1475 ( .A1(n1738), .A2(n1737), .ZN(n2019) );
  NAND2_X1 U1476 ( .A1(n1997), .A2(n1996), .ZN(n1737) );
  NAND2_X1 U1477 ( .A1(n2004), .A2(n2003), .ZN(n2011) );
  NAND2_X1 U1478 ( .A1(n1933), .A2(n1932), .ZN(n1941) );
  NAND2_X1 U1479 ( .A1(n1931), .A2(n1930), .ZN(n1932) );
  NAND2_X1 U1480 ( .A1(n1929), .A2(n1928), .ZN(n1933) );
  OR2_X1 U1481 ( .A1(n1930), .A2(n1931), .ZN(n1928) );
  XNOR2_X1 U1482 ( .A(n1929), .B(n1849), .ZN(n1856) );
  XNOR2_X1 U1483 ( .A(n1930), .B(n1931), .ZN(n1849) );
  NAND2_X1 U1484 ( .A1(n1773), .A2(n1772), .ZN(n1824) );
  NAND2_X1 U1485 ( .A1(n1813), .A2(n1812), .ZN(n1772) );
  NAND2_X1 U1486 ( .A1(n1815), .A2(n1771), .ZN(n1773) );
  OR2_X1 U1487 ( .A1(n1813), .A2(n1812), .ZN(n1771) );
  XNOR2_X1 U1488 ( .A(n1790), .B(n1789), .ZN(n1808) );
  XNOR2_X1 U1489 ( .A(n1788), .B(n1787), .ZN(n1789) );
  NOR2_X1 U1490 ( .A1(xmem_addr[4]), .A2(n2931), .ZN(n3112) );
  NAND2_X1 U1491 ( .A1(s_ready_x), .A2(s_valid_x), .ZN(n2931) );
  XNOR2_X1 U1492 ( .A(n1477), .B(n1476), .ZN(n1538) );
  NAND2_X1 U1493 ( .A1(n1808), .A2(n1807), .ZN(n2179) );
  BUF_X1 U1494 ( .A(n2831), .Z(n2575) );
  AND2_X1 U1495 ( .A1(n2908), .A2(n2817), .ZN(n3254) );
  NAND2_X1 U1496 ( .A1(n2932), .A2(n3112), .ZN(n2999) );
  INV_X1 U1497 ( .A(n2931), .ZN(n2908) );
  NAND2_X1 U1498 ( .A1(n2293), .A2(n2292), .ZN(n2391) );
  AOI21_X1 U1499 ( .B1(n2291), .B2(n2320), .A(n2290), .ZN(n2292) );
  NAND2_X1 U1500 ( .A1(n2289), .A2(n2288), .ZN(n2293) );
  CLKBUF_X1 U1501 ( .A(n2367), .Z(n2372) );
  INV_X1 U1502 ( .A(n2172), .ZN(n2173) );
  INV_X1 U1503 ( .A(n2348), .ZN(n2167) );
  INV_X1 U1504 ( .A(n2185), .ZN(n2170) );
  AOI21_X1 U1505 ( .B1(n2073), .B2(n2072), .A(n1821), .ZN(n2358) );
  AND2_X1 U1506 ( .A1(n2637), .A2(n2634), .ZN(n2652) );
  OR2_X1 U1507 ( .A1(\mac_unit_inst/adder_reg [13]), .A2(
        \mac_unit_inst/x_mult_f_reg [13]), .ZN(n2753) );
  OR2_X1 U1508 ( .A1(\mac_unit_inst/adder_reg [12]), .A2(
        \mac_unit_inst/x_mult_f_reg [12]), .ZN(n2750) );
  OR2_X1 U1509 ( .A1(n3307), .A2(n2618), .ZN(n2785) );
  CLKBUF_X1 U1510 ( .A(n2793), .Z(n2797) );
  OAI21_X1 U1511 ( .B1(n2338), .B2(n2342), .A(n2339), .ZN(n1341) );
  NAND2_X1 U1512 ( .A1(n1923), .A2(n1922), .ZN(n1876) );
  NAND2_X1 U1513 ( .A1(n1672), .A2(n1671), .ZN(n1342) );
  XNOR2_X1 U1514 ( .A(n2093), .B(n1529), .ZN(n1343) );
  NOR2_X1 U1515 ( .A1(n2027), .A2(n2026), .ZN(n1344) );
  NOR2_X1 U1516 ( .A1(n2027), .A2(n2026), .ZN(n2376) );
  XNOR2_X1 U1517 ( .A(n1352), .B(n1345), .ZN(n1791) );
  NOR2_X2 U1518 ( .A1(n3184), .A2(n2195), .ZN(n2442) );
  NOR2_X2 U1519 ( .A1(n3334), .A2(n3137), .ZN(n3230) );
  NOR2_X2 U1520 ( .A1(n3137), .A2(n3089), .ZN(n3045) );
  NOR2_X2 U1521 ( .A1(n3160), .A2(n3089), .ZN(n3067) );
  NOR2_X2 U1522 ( .A1(n3184), .A2(n3089), .ZN(n3090) );
  NOR2_X2 U1523 ( .A1(n3184), .A2(n3334), .ZN(n2447) );
  NOR2_X2 U1524 ( .A1(n3114), .A2(n2195), .ZN(n2415) );
  NOR2_X2 U1525 ( .A1(n3137), .A2(n2195), .ZN(n2457) );
  NOR2_X2 U1526 ( .A1(n3114), .A2(n3089), .ZN(n3042) );
  NOR2_X2 U1527 ( .A1(n3137), .A2(n3183), .ZN(n3157) );
  NOR2_X2 U1528 ( .A1(n3160), .A2(n3183), .ZN(n3180) );
  NOR2_X2 U1529 ( .A1(n3184), .A2(n3183), .ZN(n3204) );
  BUF_X2 U1530 ( .A(xmem_data[3]), .Z(n1869) );
  XOR2_X1 U1531 ( .A(n2129), .B(n2128), .Z(n1353) );
  XOR2_X1 U1532 ( .A(n2119), .B(n2118), .Z(n1354) );
  NOR2_X1 U1533 ( .A1(n2123), .A2(n2122), .ZN(n1355) );
  NOR2_X1 U1534 ( .A1(n2114), .A2(n2113), .ZN(n1356) );
  OR2_X1 U1535 ( .A1(n2800), .A2(n3382), .ZN(n1357) );
  OR2_X1 U1536 ( .A1(n2800), .A2(n3385), .ZN(n1358) );
  OR2_X1 U1537 ( .A1(n2800), .A2(n3381), .ZN(n1359) );
  OR2_X1 U1538 ( .A1(n2800), .A2(n3383), .ZN(n1360) );
  OR2_X1 U1539 ( .A1(n2800), .A2(n3384), .ZN(n1361) );
  OR2_X1 U1540 ( .A1(n2800), .A2(n3387), .ZN(n1362) );
  OR2_X1 U1541 ( .A1(n2800), .A2(n3378), .ZN(n1363) );
  OR2_X1 U1542 ( .A1(n2800), .A2(n3379), .ZN(n1364) );
  OR2_X1 U1543 ( .A1(n2800), .A2(n3380), .ZN(n1365) );
  OR2_X1 U1544 ( .A1(n2800), .A2(n3375), .ZN(n1366) );
  OR2_X1 U1545 ( .A1(n2800), .A2(n3386), .ZN(n1367) );
  OR2_X1 U1546 ( .A1(n2800), .A2(n3370), .ZN(n1368) );
  OR2_X1 U1547 ( .A1(n2800), .A2(n3371), .ZN(n1369) );
  OR2_X1 U1548 ( .A1(n2800), .A2(n3374), .ZN(n1370) );
  OR2_X1 U1549 ( .A1(n2800), .A2(n3372), .ZN(n1371) );
  OR2_X1 U1550 ( .A1(n2800), .A2(n3373), .ZN(n1372) );
  OR2_X1 U1551 ( .A1(n2800), .A2(n3376), .ZN(n1373) );
  OR2_X1 U1552 ( .A1(n2800), .A2(n3377), .ZN(n1374) );
  OR2_X1 U1553 ( .A1(n2800), .A2(n3388), .ZN(n1375) );
  OR2_X1 U1554 ( .A1(n1740), .A2(n1739), .ZN(n1376) );
  OR2_X1 U1555 ( .A1(n2002), .A2(n2001), .ZN(n1377) );
  NOR3_X1 U1556 ( .A1(n2221), .A2(n2220), .A3(n2219), .ZN(n1378) );
  NOR3_X1 U1557 ( .A1(n2234), .A2(n2233), .A3(n2232), .ZN(n1379) );
  NOR3_X1 U1558 ( .A1(n2247), .A2(n2246), .A3(n2245), .ZN(n1380) );
  NOR3_X1 U1559 ( .A1(n2260), .A2(n2259), .A3(n2258), .ZN(n1381) );
  NOR3_X1 U1560 ( .A1(n2273), .A2(n2272), .A3(n2271), .ZN(n1382) );
  OR2_X1 U1561 ( .A1(n1453), .A2(n1452), .ZN(n1383) );
  NOR3_X1 U1562 ( .A1(n2286), .A2(n2285), .A3(n2284), .ZN(n1384) );
  XNOR2_X1 U1563 ( .A(n2123), .B(n2122), .ZN(n1385) );
  OR2_X1 U1564 ( .A1(n2058), .A2(n2057), .ZN(n1386) );
  XNOR2_X1 U1571 ( .A(n3322), .B(n3323), .ZN(n1387) );
  XNOR2_X1 U1572 ( .A(n3391), .B(xmem_data[10]), .ZN(n1424) );
  NAND2_X2 U1573 ( .A1(n1387), .A2(n1424), .ZN(n1914) );
  INV_X2 U1574 ( .A(n3391), .ZN(n1728) );
  XNOR2_X1 U1575 ( .A(n1728), .B(fmem_data[9]), .ZN(n1411) );
  INV_X1 U1576 ( .A(n1387), .ZN(n1868) );
  INV_X2 U1577 ( .A(n1868), .ZN(n1912) );
  XNOR2_X1 U1578 ( .A(n1728), .B(fmem_data[19]), .ZN(n1425) );
  OAI22_X1 U1579 ( .A1(n1914), .A2(n1411), .B1(n1912), .B2(n1425), .ZN(n1421)
         );
  XNOR2_X1 U1580 ( .A(n3318), .B(n3315), .ZN(n1388) );
  XOR2_X1 U1581 ( .A(\DP_OP_485J1_122_4413/n1656 ), .B(xmem_data[16]), .Z(
        n1389) );
  OR2_X2 U1582 ( .A1(n1388), .A2(n1389), .ZN(n1581) );
  BUF_X2 U1583 ( .A(\DP_OP_485J1_122_4413/n1655 ), .Z(n1579) );
  XNOR2_X1 U1584 ( .A(n1579), .B(fmem_data[3]), .ZN(n1392) );
  XNOR2_X1 U1585 ( .A(n1579), .B(fmem_data[4]), .ZN(n1416) );
  OAI22_X1 U1586 ( .A1(n1581), .A2(n1392), .B1(n1546), .B2(n1416), .ZN(n1420)
         );
  XNOR2_X1 U1587 ( .A(\DP_OP_485J1_122_4413/n1656 ), .B(xmem_data[14]), .ZN(
        n1390) );
  XNOR2_X1 U1588 ( .A(\DP_OP_485J1_122_4413/n1657 ), .B(n3316), .ZN(n1391) );
  OR2_X2 U1589 ( .A1(n1390), .A2(n1391), .ZN(n1577) );
  BUF_X2 U1590 ( .A(\DP_OP_485J1_122_4413/n1656 ), .Z(n1557) );
  XNOR2_X1 U1591 ( .A(n1557), .B(fmem_data[5]), .ZN(n1397) );
  XNOR2_X1 U1592 ( .A(n1557), .B(fmem_data[6]), .ZN(n1417) );
  OAI22_X1 U1593 ( .A1(n1577), .A2(n1397), .B1(n1629), .B2(n1417), .ZN(n1419)
         );
  XNOR2_X1 U1594 ( .A(n1579), .B(fmem_data[2]), .ZN(n1403) );
  OAI22_X1 U1595 ( .A1(n1581), .A2(n1403), .B1(n1546), .B2(n1392), .ZN(n1434)
         );
  XNOR2_X1 U1596 ( .A(xmem_data[19]), .B(n3324), .ZN(n1393) );
  XNOR2_X1 U1597 ( .A(xmem_data[18]), .B(\DP_OP_485J1_122_4413/n1655 ), .ZN(
        n1394) );
  NAND2_X2 U1598 ( .A1(n1393), .A2(n1394), .ZN(n1613) );
  XNOR2_X1 U1599 ( .A(\DP_OP_485J1_122_4413/n1204 ), .B(n1607), .ZN(n1396) );
  INV_X1 U1600 ( .A(n1394), .ZN(n1395) );
  INV_X2 U1601 ( .A(n1395), .ZN(n1614) );
  XNOR2_X1 U1602 ( .A(xmem_data[19]), .B(fmem_data[1]), .ZN(n1409) );
  OAI22_X1 U1603 ( .A1(n1613), .A2(n1396), .B1(n1614), .B2(n1409), .ZN(n1433)
         );
  XNOR2_X1 U1604 ( .A(n1557), .B(fmem_data[4]), .ZN(n1404) );
  OAI22_X1 U1605 ( .A1(n1577), .A2(n1404), .B1(n1629), .B2(n1397), .ZN(n1432)
         );
  INV_X1 U1606 ( .A(n3319), .ZN(n1398) );
  XOR2_X1 U1607 ( .A(\DP_OP_485J1_122_4413/n1657 ), .B(n1398), .Z(n1651) );
  XNOR2_X2 U1608 ( .A(n3320), .B(xmem_data[12]), .ZN(n1653) );
  NAND2_X1 U1609 ( .A1(n1651), .A2(n1653), .ZN(n1646) );
  BUF_X1 U1610 ( .A(n1646), .Z(n1438) );
  INV_X2 U1611 ( .A(n3327), .ZN(n1649) );
  XNOR2_X1 U1612 ( .A(n1649), .B(fmem_data[6]), .ZN(n1437) );
  XNOR2_X1 U1613 ( .A(n1649), .B(fmem_data[7]), .ZN(n1410) );
  OR2_X1 U1614 ( .A1(n1410), .A2(n1653), .ZN(n1402) );
  OAI21_X1 U1615 ( .B1(n1438), .B2(n1437), .A(n1402), .ZN(n1401) );
  XNOR2_X1 U1616 ( .A(xmem_data[7]), .B(xmem_data[8]), .ZN(n1400) );
  XOR2_X1 U1617 ( .A(xmem_data[9]), .B(xmem_data[8]), .Z(n1399) );
  NAND2_X1 U1618 ( .A1(n1400), .A2(n1399), .ZN(n1702) );
  BUF_X2 U1619 ( .A(n1702), .Z(n1893) );
  XNOR2_X1 U1620 ( .A(n1837), .B(fmem_data[9]), .ZN(n1465) );
  BUF_X2 U1621 ( .A(n1400), .Z(n1891) );
  XNOR2_X1 U1622 ( .A(n1837), .B(fmem_data[19]), .ZN(n1414) );
  OAI22_X1 U1623 ( .A1(n1893), .A2(n1465), .B1(n1891), .B2(n1414), .ZN(n1436)
         );
  AND2_X1 U1624 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1395), .ZN(n1435) );
  OR2_X1 U1625 ( .A1(n1436), .A2(n1435), .ZN(n1474) );
  NAND2_X1 U1626 ( .A1(n1401), .A2(n1474), .ZN(n1406) );
  OAI21_X1 U1627 ( .B1(n1438), .B2(n1437), .A(n1402), .ZN(n1475) );
  XNOR2_X1 U1628 ( .A(n1579), .B(fmem_data[1]), .ZN(n1440) );
  OAI22_X1 U1629 ( .A1(n1581), .A2(n1440), .B1(n1546), .B2(n1403), .ZN(n1462)
         );
  XNOR2_X1 U1630 ( .A(n1557), .B(fmem_data[3]), .ZN(n1463) );
  OAI22_X1 U1631 ( .A1(n1577), .A2(n1463), .B1(n1629), .B2(n1404), .ZN(n1461)
         );
  XNOR2_X1 U1632 ( .A(n1728), .B(fmem_data[7]), .ZN(n1459) );
  XNOR2_X1 U1633 ( .A(n1728), .B(fmem_data[8]), .ZN(n1412) );
  OAI22_X1 U1634 ( .A1(n1914), .A2(n1459), .B1(n1912), .B2(n1412), .ZN(n1460)
         );
  OAI21_X1 U1635 ( .B1(n1475), .B2(n1474), .A(n1476), .ZN(n1405) );
  NAND2_X1 U1636 ( .A1(n1406), .A2(n1405), .ZN(n1454) );
  NAND2_X1 U1637 ( .A1(n1383), .A2(n1454), .ZN(n1408) );
  NAND2_X1 U1638 ( .A1(n1408), .A2(n1407), .ZN(n1528) );
  XNOR2_X1 U1639 ( .A(xmem_data[19]), .B(fmem_data[2]), .ZN(n1418) );
  OAI22_X1 U1640 ( .A1(n1613), .A2(n1409), .B1(n1614), .B2(n1418), .ZN(n1512)
         );
  INV_X1 U1641 ( .A(n1512), .ZN(n1451) );
  XNOR2_X1 U1642 ( .A(n1649), .B(fmem_data[8]), .ZN(n1423) );
  OAI22_X1 U1643 ( .A1(n1438), .A2(n1410), .B1(n1653), .B2(n1423), .ZN(n1450)
         );
  OAI22_X1 U1644 ( .A1(n1914), .A2(n1412), .B1(n1912), .B2(n1411), .ZN(n1431)
         );
  OR2_X1 U1645 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n3326), .ZN(n1413) );
  OAI22_X1 U1646 ( .A1(n1613), .A2(n3326), .B1(n1413), .B2(n1614), .ZN(n1430)
         );
  AOI21_X1 U1647 ( .B1(n1831), .B2(n1891), .A(n1414), .ZN(n1415) );
  INV_X1 U1648 ( .A(n1415), .ZN(n1429) );
  XNOR2_X1 U1649 ( .A(n1528), .B(n1527), .ZN(n1531) );
  XNOR2_X1 U1650 ( .A(n1579), .B(fmem_data[5]), .ZN(n1518) );
  OAI22_X1 U1651 ( .A1(n1581), .A2(n1416), .B1(n1546), .B2(n1518), .ZN(n1515)
         );
  XNOR2_X1 U1652 ( .A(n1557), .B(fmem_data[7]), .ZN(n1519) );
  OAI22_X1 U1653 ( .A1(n1577), .A2(n1417), .B1(n1629), .B2(n1519), .ZN(n1514)
         );
  XNOR2_X1 U1654 ( .A(xmem_data[19]), .B(fmem_data[3]), .ZN(n1516) );
  OAI22_X1 U1655 ( .A1(n1613), .A2(n1418), .B1(n1614), .B2(n1516), .ZN(n1513)
         );
  FA_X1 U1656 ( .A(n1421), .B(n1420), .CI(n1419), .CO(n1522), .S(n1453) );
  XNOR2_X1 U1657 ( .A(n1523), .B(n1522), .ZN(n1428) );
  NAND2_X1 U1658 ( .A1(n1651), .A2(n1653), .ZN(n1634) );
  XNOR2_X1 U1659 ( .A(n1649), .B(fmem_data[9]), .ZN(n1520) );
  OR2_X1 U1660 ( .A1(n1520), .A2(n1653), .ZN(n1422) );
  OAI21_X1 U1661 ( .B1(n1634), .B2(n1423), .A(n1422), .ZN(n1511) );
  INV_X1 U1662 ( .A(n1424), .ZN(n1426) );
  AOI21_X1 U1663 ( .B1(n1426), .B2(n1912), .A(n1425), .ZN(n1427) );
  INV_X1 U1664 ( .A(n1427), .ZN(n1510) );
  XNOR2_X1 U1665 ( .A(n1428), .B(n1521), .ZN(n1530) );
  XNOR2_X1 U1666 ( .A(n1531), .B(n1530), .ZN(n2090) );
  FA_X1 U1667 ( .A(n1431), .B(n1430), .CI(n1429), .CO(n1449), .S(n1479) );
  FA_X1 U1668 ( .A(n1434), .B(n1433), .CI(n1432), .CO(n1452), .S(n1478) );
  NOR2_X1 U1669 ( .A1(n1479), .A2(n1478), .ZN(n1448) );
  XNOR2_X1 U1670 ( .A(n1436), .B(n1435), .ZN(n1484) );
  XNOR2_X1 U1671 ( .A(n1649), .B(fmem_data[5]), .ZN(n1467) );
  OAI22_X1 U1672 ( .A1(n1438), .A2(n1467), .B1(n1653), .B2(n1437), .ZN(n1483)
         );
  OR2_X1 U1673 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n3318), .ZN(n1439) );
  OAI22_X1 U1674 ( .A1(n1581), .A2(n3318), .B1(n1439), .B2(n1546), .ZN(n1490)
         );
  XNOR2_X1 U1675 ( .A(\DP_OP_485J1_122_4413/n1204 ), .B(n1579), .ZN(n1441) );
  OAI22_X1 U1676 ( .A1(n1581), .A2(n1441), .B1(n1546), .B2(n1440), .ZN(n1489)
         );
  INV_X1 U1677 ( .A(n3317), .ZN(n1442) );
  XNOR2_X1 U1678 ( .A(n1442), .B(n3321), .ZN(n1444) );
  INV_X1 U1679 ( .A(n1444), .ZN(n1885) );
  XNOR2_X1 U1680 ( .A(xmem_data[7]), .B(xmem_data[6]), .ZN(n1443) );
  OR2_X2 U1681 ( .A1(n1444), .A2(n1443), .ZN(n1887) );
  INV_X1 U1682 ( .A(n3329), .ZN(n1866) );
  XNOR2_X1 U1683 ( .A(n1866), .B(fmem_data[19]), .ZN(n1457) );
  AOI21_X1 U1684 ( .B1(n1885), .B2(n1887), .A(n1457), .ZN(n1445) );
  INV_X1 U1685 ( .A(n1445), .ZN(n1488) );
  INV_X1 U1686 ( .A(n1480), .ZN(n1447) );
  OAI21_X1 U1687 ( .B1(n1448), .B2(n1447), .A(n1446), .ZN(n1536) );
  FA_X1 U1688 ( .A(n1451), .B(n1450), .CI(n1449), .CO(n1527), .S(n1535) );
  XNOR2_X1 U1689 ( .A(n1453), .B(n1452), .ZN(n1455) );
  XNOR2_X1 U1690 ( .A(n1455), .B(n1454), .ZN(n1534) );
  INV_X1 U1691 ( .A(n2089), .ZN(n1456) );
  XNOR2_X1 U1692 ( .A(n2090), .B(n1456), .ZN(n2039) );
  BUF_X1 U1693 ( .A(xmem_data[7]), .Z(n1745) );
  XNOR2_X1 U1694 ( .A(n1745), .B(fmem_data[9]), .ZN(n1624) );
  OAI22_X1 U1695 ( .A1(n1887), .A2(n1624), .B1(n1885), .B2(n1457), .ZN(n1492)
         );
  INV_X1 U1696 ( .A(n1546), .ZN(n1458) );
  AND2_X1 U1697 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1458), .ZN(n1491) );
  OR2_X1 U1698 ( .A1(n1492), .A2(n1491), .ZN(n1637) );
  XNOR2_X1 U1699 ( .A(n1728), .B(fmem_data[6]), .ZN(n1493) );
  OAI22_X1 U1700 ( .A1(n1914), .A2(n1493), .B1(n1912), .B2(n1459), .ZN(n1636)
         );
  XNOR2_X1 U1701 ( .A(n1557), .B(fmem_data[1]), .ZN(n1497) );
  XNOR2_X1 U1702 ( .A(n1557), .B(fmem_data[2]), .ZN(n1464) );
  OAI22_X1 U1703 ( .A1(n1577), .A2(n1497), .B1(n1629), .B2(n1464), .ZN(n1622)
         );
  XNOR2_X1 U1704 ( .A(n1837), .B(fmem_data[7]), .ZN(n1630) );
  XNOR2_X1 U1705 ( .A(n1837), .B(fmem_data[8]), .ZN(n1466) );
  OAI22_X1 U1706 ( .A1(n1893), .A2(n1630), .B1(n1891), .B2(n1466), .ZN(n1621)
         );
  NAND2_X1 U1707 ( .A1(n1651), .A2(n1653), .ZN(n1549) );
  XNOR2_X1 U1708 ( .A(n1649), .B(fmem_data[3]), .ZN(n1625) );
  XNOR2_X1 U1709 ( .A(n1649), .B(fmem_data[4]), .ZN(n1468) );
  OAI22_X1 U1710 ( .A1(n1549), .A2(n1625), .B1(n1653), .B2(n1468), .ZN(n1620)
         );
  FA_X1 U1711 ( .A(n1462), .B(n1461), .CI(n1460), .CO(n1476), .S(n1505) );
  INV_X1 U1712 ( .A(n1505), .ZN(n1470) );
  OAI22_X1 U1713 ( .A1(n1577), .A2(n1464), .B1(n1629), .B2(n1463), .ZN(n1487)
         );
  OAI22_X1 U1714 ( .A1(n1831), .A2(n1466), .B1(n1891), .B2(n1465), .ZN(n1486)
         );
  OAI22_X1 U1715 ( .A1(n1549), .A2(n1468), .B1(n1653), .B2(n1467), .ZN(n1485)
         );
  INV_X1 U1716 ( .A(n1504), .ZN(n1469) );
  NAND2_X1 U1717 ( .A1(n1470), .A2(n1469), .ZN(n1471) );
  NAND2_X1 U1718 ( .A1(n1507), .A2(n1471), .ZN(n1473) );
  NAND2_X1 U1719 ( .A1(n1505), .A2(n1504), .ZN(n1472) );
  NAND2_X1 U1720 ( .A1(n1473), .A2(n1472), .ZN(n1539) );
  XNOR2_X1 U1721 ( .A(n1479), .B(n1478), .ZN(n1481) );
  XNOR2_X1 U1722 ( .A(n1481), .B(n1480), .ZN(n1537) );
  INV_X1 U1723 ( .A(n1533), .ZN(n2077) );
  FA_X1 U1724 ( .A(n1484), .B(n1483), .CI(n1482), .CO(n1480), .S(n1680) );
  FA_X1 U1725 ( .A(n1487), .B(n1486), .CI(n1485), .CO(n1504), .S(n1640) );
  FA_X1 U1726 ( .A(n1490), .B(n1489), .CI(n1488), .CO(n1482), .S(n1638) );
  XNOR2_X1 U1727 ( .A(n1492), .B(n1491), .ZN(n1675) );
  XNOR2_X1 U1728 ( .A(n1728), .B(fmem_data[5]), .ZN(n1623) );
  OAI22_X1 U1729 ( .A1(n1914), .A2(n1623), .B1(n1912), .B2(n1493), .ZN(n1674)
         );
  INV_X1 U1730 ( .A(xmem_data[5]), .ZN(n1494) );
  XNOR2_X1 U1731 ( .A(xmem_data[4]), .B(n1494), .ZN(n1627) );
  INV_X1 U1732 ( .A(n1627), .ZN(n1495) );
  XNOR2_X1 U1733 ( .A(xmem_data[4]), .B(xmem_data[3]), .ZN(n1626) );
  BUF_X2 U1734 ( .A(xmem_data[5]), .Z(n1894) );
  XNOR2_X1 U1735 ( .A(n1894), .B(fmem_data[19]), .ZN(n1628) );
  AOI21_X1 U1736 ( .B1(n1495), .B2(n1909), .A(n1628), .ZN(n1496) );
  INV_X1 U1737 ( .A(n1496), .ZN(n1666) );
  XNOR2_X1 U1738 ( .A(\DP_OP_485J1_122_4413/n1204 ), .B(n1557), .ZN(n1498) );
  OAI22_X1 U1739 ( .A1(n1498), .A2(n1577), .B1(n1629), .B2(n1497), .ZN(n1667)
         );
  OR2_X1 U1740 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1351), .ZN(n1499) );
  OAI22_X1 U1741 ( .A1(n1577), .A2(n1351), .B1(n1499), .B2(n1629), .ZN(n1669)
         );
  OAI21_X1 U1742 ( .B1(n1666), .B2(n1667), .A(n1669), .ZN(n1501) );
  NAND2_X1 U1743 ( .A1(n1666), .A2(n1667), .ZN(n1500) );
  NAND2_X1 U1744 ( .A1(n1501), .A2(n1500), .ZN(n1673) );
  OAI21_X1 U1745 ( .B1(n1640), .B2(n1638), .A(n1639), .ZN(n1503) );
  NAND2_X1 U1746 ( .A1(n1640), .A2(n1638), .ZN(n1502) );
  NAND2_X1 U1747 ( .A1(n1503), .A2(n1502), .ZN(n1679) );
  XNOR2_X1 U1748 ( .A(n1505), .B(n1504), .ZN(n1506) );
  XNOR2_X1 U1749 ( .A(n1507), .B(n1506), .ZN(n1681) );
  OAI21_X1 U1750 ( .B1(n1680), .B2(n1679), .A(n1681), .ZN(n1509) );
  NAND2_X1 U1751 ( .A1(n1679), .A2(n1680), .ZN(n1508) );
  AND2_X2 U1752 ( .A1(n1509), .A2(n1508), .ZN(n2786) );
  NOR2_X1 U1753 ( .A1(n2077), .A2(n2786), .ZN(n2038) );
  FA_X1 U1754 ( .A(n1512), .B(n1511), .CI(n1510), .CO(n1543), .S(n1521) );
  FA_X1 U1755 ( .A(n1515), .B(n1514), .CI(n1513), .CO(n1541), .S(n1523) );
  XNOR2_X1 U1756 ( .A(xmem_data[19]), .B(fmem_data[4]), .ZN(n1552) );
  OAI22_X1 U1757 ( .A1(n1613), .A2(n1516), .B1(n1614), .B2(n1552), .ZN(n1561)
         );
  INV_X1 U1758 ( .A(n1561), .ZN(n1542) );
  XNOR2_X1 U1759 ( .A(n1541), .B(n1542), .ZN(n1517) );
  XNOR2_X1 U1760 ( .A(n1543), .B(n1517), .ZN(n1571) );
  XNOR2_X1 U1761 ( .A(n1579), .B(fmem_data[6]), .ZN(n1547) );
  OAI22_X1 U1762 ( .A1(n1581), .A2(n1518), .B1(n1546), .B2(n1547), .ZN(n1555)
         );
  XNOR2_X1 U1763 ( .A(n1557), .B(fmem_data[8]), .ZN(n1551) );
  OAI22_X1 U1764 ( .A1(n1577), .A2(n1519), .B1(n1629), .B2(n1551), .ZN(n1554)
         );
  XNOR2_X1 U1765 ( .A(n1649), .B(fmem_data[19]), .ZN(n1548) );
  OAI22_X1 U1766 ( .A1(n1634), .A2(n1520), .B1(n1653), .B2(n1548), .ZN(n1553)
         );
  INV_X1 U1767 ( .A(n1521), .ZN(n1525) );
  OAI21_X1 U1768 ( .B1(n1526), .B2(n1525), .A(n1524), .ZN(n1569) );
  OAI21_X1 U1769 ( .B1(n1528), .B2(n1527), .A(n1530), .ZN(n1594) );
  NAND2_X1 U1770 ( .A1(n1528), .A2(n1527), .ZN(n1593) );
  AND2_X1 U1771 ( .A1(n1594), .A2(n1593), .ZN(n1529) );
  XNOR2_X1 U1772 ( .A(n2093), .B(n1529), .ZN(n2040) );
  XNOR2_X1 U1773 ( .A(n1531), .B(n1530), .ZN(n2076) );
  AND2_X1 U1774 ( .A1(n2076), .A2(n2089), .ZN(n2041) );
  OAI22_X1 U1775 ( .A1(n2039), .A2(n2038), .B1(n2040), .B2(n2041), .ZN(n1532)
         );
  INV_X1 U1776 ( .A(n1532), .ZN(n2047) );
  XNOR2_X1 U1777 ( .A(n2786), .B(n1533), .ZN(n2035) );
  FA_X1 U1778 ( .A(n1536), .B(n1535), .CI(n1534), .CO(n2089), .S(n2080) );
  NOR2_X1 U1779 ( .A1(n2035), .A2(n2080), .ZN(n2037) );
  FA_X1 U1780 ( .A(n1539), .B(n1538), .CI(n1537), .CO(n1533), .S(n2788) );
  NOR2_X1 U1781 ( .A1(n2788), .A2(n2786), .ZN(n2143) );
  NOR2_X1 U1782 ( .A1(n2037), .A2(n2143), .ZN(n1540) );
  NAND2_X1 U1783 ( .A1(n2047), .A2(n1540), .ZN(n1619) );
  OAI21_X1 U1784 ( .B1(n1543), .B2(n1542), .A(n1541), .ZN(n1545) );
  NAND2_X1 U1785 ( .A1(n1543), .A2(n1542), .ZN(n1544) );
  NAND2_X1 U1786 ( .A1(n1545), .A2(n1544), .ZN(n1568) );
  XNOR2_X1 U1787 ( .A(n1579), .B(fmem_data[7]), .ZN(n1556) );
  OAI22_X1 U1788 ( .A1(n1581), .A2(n1547), .B1(n1601), .B2(n1556), .ZN(n1562)
         );
  AOI21_X1 U1789 ( .B1(n1549), .B2(n1653), .A(n1548), .ZN(n1550) );
  INV_X1 U1790 ( .A(n1550), .ZN(n1560) );
  XNOR2_X1 U1791 ( .A(n1557), .B(fmem_data[9]), .ZN(n1558) );
  OAI22_X1 U1792 ( .A1(n1577), .A2(n1551), .B1(n1629), .B2(n1558), .ZN(n1565)
         );
  XNOR2_X1 U1793 ( .A(xmem_data[19]), .B(fmem_data[5]), .ZN(n1559) );
  OAI22_X1 U1794 ( .A1(n1613), .A2(n1552), .B1(n1614), .B2(n1559), .ZN(n1564)
         );
  FA_X1 U1795 ( .A(n1555), .B(n1554), .CI(n1553), .CO(n1563), .S(n1570) );
  XNOR2_X1 U1796 ( .A(n1579), .B(fmem_data[8]), .ZN(n1580) );
  OAI22_X1 U1797 ( .A1(n1581), .A2(n1556), .B1(n1601), .B2(n1580), .ZN(n1574)
         );
  XNOR2_X1 U1798 ( .A(n1557), .B(fmem_data[19]), .ZN(n1576) );
  OAI22_X1 U1799 ( .A1(n1577), .A2(n1558), .B1(n1629), .B2(n1576), .ZN(n1573)
         );
  XNOR2_X1 U1800 ( .A(xmem_data[19]), .B(fmem_data[6]), .ZN(n1575) );
  OAI22_X1 U1801 ( .A1(n1613), .A2(n1559), .B1(n1614), .B2(n1575), .ZN(n1588)
         );
  INV_X1 U1802 ( .A(n1588), .ZN(n1572) );
  FA_X1 U1803 ( .A(n1562), .B(n1561), .CI(n1560), .CO(n1583), .S(n1567) );
  FA_X1 U1804 ( .A(n1565), .B(n1564), .CI(n1563), .CO(n1582), .S(n1566) );
  FA_X1 U1805 ( .A(n1568), .B(n1567), .CI(n1566), .CO(n2097), .S(n2096) );
  FA_X1 U1806 ( .A(n1571), .B(n1570), .CI(n1569), .CO(n2095), .S(n2093) );
  FA_X1 U1807 ( .A(n1574), .B(n1573), .CI(n1572), .CO(n1592), .S(n1584) );
  XNOR2_X1 U1808 ( .A(n1607), .B(fmem_data[7]), .ZN(n1585) );
  OAI22_X1 U1809 ( .A1(n1613), .A2(n1575), .B1(n1614), .B2(n1585), .ZN(n1591)
         );
  AOI21_X1 U1810 ( .B1(n1577), .B2(n1629), .A(n1576), .ZN(n1578) );
  INV_X1 U1811 ( .A(n1578), .ZN(n1589) );
  XNOR2_X1 U1812 ( .A(n1579), .B(fmem_data[9]), .ZN(n1586) );
  OAI22_X1 U1813 ( .A1(n1581), .A2(n1580), .B1(n1601), .B2(n1586), .ZN(n1587)
         );
  FA_X1 U1814 ( .A(n1584), .B(n1583), .CI(n1582), .CO(n2113), .S(n2098) );
  XOR2_X1 U1815 ( .A(n2114), .B(n2113), .Z(n2054) );
  XNOR2_X1 U1816 ( .A(n1607), .B(fmem_data[8]), .ZN(n1599) );
  OAI22_X1 U1817 ( .A1(n1613), .A2(n1585), .B1(n1614), .B2(n1599), .ZN(n1605)
         );
  INV_X1 U1818 ( .A(n1605), .ZN(n1598) );
  XNOR2_X1 U1819 ( .A(n1579), .B(fmem_data[19]), .ZN(n1600) );
  OAI22_X1 U1820 ( .A1(n1581), .A2(n1586), .B1(n1601), .B2(n1600), .ZN(n1597)
         );
  FA_X1 U1821 ( .A(n1589), .B(n1588), .CI(n1587), .CO(n1596), .S(n1590) );
  FA_X1 U1822 ( .A(n1592), .B(n1591), .CI(n1590), .CO(n2118), .S(n2114) );
  HA_X1 U1823 ( .A(n2119), .B(n2118), .S(n2056) );
  AND2_X1 U1824 ( .A1(n2054), .A2(n2056), .ZN(n2052) );
  OAI21_X1 U1825 ( .B1(n2050), .B2(n2051), .A(n2052), .ZN(n2060) );
  HA_X1 U1826 ( .A(n2096), .B(n2095), .CO(n2051), .S(n2049) );
  NAND2_X1 U1827 ( .A1(n1594), .A2(n1593), .ZN(n2092) );
  AND2_X1 U1828 ( .A1(n2093), .A2(n2092), .ZN(n2048) );
  NOR2_X1 U1829 ( .A1(n2049), .A2(n2048), .ZN(n1595) );
  NOR2_X1 U1830 ( .A1(n1595), .A2(n2060), .ZN(n1618) );
  FA_X1 U1831 ( .A(n1598), .B(n1597), .CI(n1596), .CO(n2121), .S(n2119) );
  XNOR2_X1 U1832 ( .A(n1607), .B(fmem_data[9]), .ZN(n1608) );
  OAI22_X1 U1833 ( .A1(n1613), .A2(n1599), .B1(n1614), .B2(n1608), .ZN(n1606)
         );
  AOI21_X1 U1834 ( .B1(n1601), .B2(n1581), .A(n1600), .ZN(n1602) );
  INV_X1 U1835 ( .A(n1602), .ZN(n1604) );
  HA_X1 U1836 ( .A(n2121), .B(n2120), .S(n1603) );
  INV_X1 U1837 ( .A(n1603), .ZN(n1611) );
  FA_X1 U1838 ( .A(n1606), .B(n1605), .CI(n1604), .CO(n2123), .S(n2120) );
  XNOR2_X1 U1839 ( .A(n1607), .B(fmem_data[19]), .ZN(n1612) );
  OAI22_X1 U1840 ( .A1(n1613), .A2(n1608), .B1(n1614), .B2(n1612), .ZN(n2128)
         );
  INV_X1 U1841 ( .A(n2128), .ZN(n2122) );
  HA_X1 U1842 ( .A(n2123), .B(n2122), .S(n1609) );
  INV_X1 U1843 ( .A(n1609), .ZN(n1610) );
  NOR2_X1 U1844 ( .A1(n1611), .A2(n1610), .ZN(n1617) );
  AOI21_X1 U1845 ( .B1(n1614), .B2(n1613), .A(n1612), .ZN(n1615) );
  INV_X1 U1846 ( .A(n1615), .ZN(n2129) );
  NAND2_X1 U1847 ( .A1(n1618), .A2(n2063), .ZN(n2065) );
  NOR2_X1 U1848 ( .A1(n1619), .A2(n2065), .ZN(n2068) );
  FA_X1 U1849 ( .A(n1622), .B(n1621), .CI(n1620), .CO(n1635), .S(n1678) );
  XNOR2_X1 U1850 ( .A(n1728), .B(fmem_data[4]), .ZN(n1632) );
  OAI22_X1 U1851 ( .A1(n1914), .A2(n1632), .B1(n1912), .B2(n1623), .ZN(n1665)
         );
  XNOR2_X1 U1852 ( .A(n1745), .B(fmem_data[8]), .ZN(n1631) );
  OAI22_X1 U1853 ( .A1(n1887), .A2(n1631), .B1(n1885), .B2(n1624), .ZN(n1664)
         );
  XNOR2_X1 U1854 ( .A(n1649), .B(fmem_data[2]), .ZN(n1633) );
  OAI22_X1 U1855 ( .A1(n1646), .A2(n1633), .B1(n1653), .B2(n1625), .ZN(n1663)
         );
  NAND2_X1 U1856 ( .A1(n1627), .A2(n1626), .ZN(n1750) );
  BUF_X1 U1857 ( .A(n1750), .Z(n1833) );
  XNOR2_X1 U1858 ( .A(n1894), .B(fmem_data[9]), .ZN(n1694) );
  OAI22_X1 U1859 ( .A1(n1833), .A2(n1694), .B1(n1909), .B2(n1628), .ZN(n1643)
         );
  AND2_X1 U1860 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1391), .ZN(n1642) );
  OR2_X1 U1861 ( .A1(n1643), .A2(n1642), .ZN(n1710) );
  XNOR2_X1 U1862 ( .A(n1837), .B(fmem_data[6]), .ZN(n1644) );
  OAI22_X1 U1863 ( .A1(n1893), .A2(n1644), .B1(n1891), .B2(n1630), .ZN(n1709)
         );
  XNOR2_X1 U1864 ( .A(n1745), .B(fmem_data[7]), .ZN(n1700) );
  OAI22_X1 U1865 ( .A1(n1887), .A2(n1700), .B1(n1885), .B2(n1631), .ZN(n1692)
         );
  XNOR2_X1 U1866 ( .A(n1728), .B(fmem_data[3]), .ZN(n1693) );
  OAI22_X1 U1867 ( .A1(n1914), .A2(n1693), .B1(n1912), .B2(n1632), .ZN(n1691)
         );
  XNOR2_X1 U1868 ( .A(n1649), .B(fmem_data[1]), .ZN(n1647) );
  OAI22_X1 U1869 ( .A1(n1634), .A2(n1647), .B1(n1653), .B2(n1633), .ZN(n1690)
         );
  FA_X1 U1870 ( .A(n1637), .B(n1636), .CI(n1635), .CO(n1507), .S(n1684) );
  XNOR2_X1 U1871 ( .A(n1639), .B(n1638), .ZN(n1641) );
  XNOR2_X1 U1872 ( .A(n1641), .B(n1640), .ZN(n1683) );
  XNOR2_X1 U1873 ( .A(n1643), .B(n1642), .ZN(n1719) );
  XNOR2_X1 U1874 ( .A(n1837), .B(fmem_data[5]), .ZN(n1695) );
  OAI22_X1 U1875 ( .A1(n1831), .A2(n1695), .B1(n1891), .B2(n1644), .ZN(n1718)
         );
  XNOR2_X1 U1876 ( .A(\DP_OP_485J1_122_4413/n1204 ), .B(n1649), .ZN(n1645) );
  NOR2_X1 U1877 ( .A1(n1646), .A2(n1645), .ZN(n1660) );
  OR2_X1 U1878 ( .A1(n1647), .A2(n1653), .ZN(n1656) );
  INV_X1 U1879 ( .A(n1656), .ZN(n1648) );
  NOR2_X1 U1880 ( .A1(n1660), .A2(n1648), .ZN(n1723) );
  INV_X1 U1881 ( .A(n1653), .ZN(n1699) );
  NOR2_X1 U1882 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n3327), .ZN(n1650) );
  NAND2_X1 U1883 ( .A1(n1699), .A2(n1650), .ZN(n1657) );
  INV_X1 U1884 ( .A(n1651), .ZN(n1652) );
  NOR2_X1 U1885 ( .A1(n1652), .A2(n3327), .ZN(n1654) );
  NAND2_X1 U1886 ( .A1(n1654), .A2(n1653), .ZN(n1655) );
  NAND2_X1 U1887 ( .A1(n1657), .A2(n1655), .ZN(n1721) );
  INV_X1 U1888 ( .A(n1721), .ZN(n1662) );
  NAND3_X1 U1889 ( .A1(n1657), .A2(n1656), .A3(n1655), .ZN(n1659) );
  XNOR2_X1 U1890 ( .A(n1869), .B(fmem_data[19]), .ZN(n1696) );
  AOI21_X1 U1891 ( .B1(n1791), .B2(n1882), .A(n1696), .ZN(n1720) );
  INV_X1 U1892 ( .A(n1720), .ZN(n1658) );
  OAI21_X1 U1893 ( .B1(n1660), .B2(n1659), .A(n1658), .ZN(n1661) );
  OAI21_X1 U1894 ( .B1(n1723), .B2(n1662), .A(n1661), .ZN(n1717) );
  FA_X1 U1895 ( .A(n1665), .B(n1664), .CI(n1663), .CO(n1677), .S(n1687) );
  XNOR2_X1 U1896 ( .A(n1667), .B(n1666), .ZN(n1668) );
  XNOR2_X1 U1897 ( .A(n1669), .B(n1668), .ZN(n1686) );
  OR2_X1 U1898 ( .A1(n1687), .A2(n1686), .ZN(n1670) );
  NAND2_X1 U1899 ( .A1(n1689), .A2(n1670), .ZN(n1672) );
  NAND2_X1 U1900 ( .A1(n1672), .A2(n1671), .ZN(n2023) );
  FA_X1 U1901 ( .A(n1675), .B(n1674), .CI(n1673), .CO(n1639), .S(n2022) );
  FA_X1 U1902 ( .A(n1678), .B(n1677), .CI(n1676), .CO(n1685), .S(n2021) );
  XNOR2_X1 U1903 ( .A(n1680), .B(n1679), .ZN(n1682) );
  XNOR2_X1 U1904 ( .A(n1682), .B(n1681), .ZN(n2029) );
  FA_X1 U1905 ( .A(n1685), .B(n1684), .CI(n1683), .CO(n2028), .S(n2027) );
  NOR2_X1 U1906 ( .A1(n2029), .A2(n2028), .ZN(n2392) );
  NOR2_X1 U1907 ( .A1(n2376), .A2(n2392), .ZN(n2031) );
  FA_X1 U1908 ( .A(n2023), .B(n2022), .CI(n2021), .S(n2018) );
  FA_X1 U1909 ( .A(n1692), .B(n1691), .CI(n1690), .CO(n1708), .S(n1714) );
  XNOR2_X1 U1910 ( .A(n1728), .B(fmem_data[2]), .ZN(n1704) );
  OAI22_X1 U1911 ( .A1(n1914), .A2(n1704), .B1(n1912), .B2(n1693), .ZN(n1726)
         );
  XNOR2_X1 U1912 ( .A(n1894), .B(fmem_data[8]), .ZN(n1701) );
  OAI22_X1 U1913 ( .A1(n1833), .A2(n1701), .B1(n1909), .B2(n1694), .ZN(n1725)
         );
  XNOR2_X1 U1914 ( .A(n1837), .B(fmem_data[4]), .ZN(n1703) );
  OAI22_X1 U1915 ( .A1(n1831), .A2(n1703), .B1(n1891), .B2(n1695), .ZN(n1724)
         );
  OR2_X1 U1916 ( .A1(n1791), .A2(n1799), .ZN(n1779) );
  XNOR2_X1 U1917 ( .A(n1869), .B(fmem_data[9]), .ZN(n1883) );
  INV_X1 U1918 ( .A(n1696), .ZN(n1697) );
  NAND2_X1 U1919 ( .A1(n1799), .A2(n1697), .ZN(n1698) );
  OAI21_X1 U1920 ( .B1(n1779), .B2(n1883), .A(n1698), .ZN(n1733) );
  AND2_X1 U1921 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1699), .ZN(n1732) );
  OR2_X1 U1922 ( .A1(n1733), .A2(n1732), .ZN(n1988) );
  XNOR2_X1 U1923 ( .A(n1745), .B(fmem_data[6]), .ZN(n1731) );
  OAI22_X1 U1924 ( .A1(n1887), .A2(n1731), .B1(n1885), .B2(n1700), .ZN(n1987)
         );
  XNOR2_X1 U1925 ( .A(n1894), .B(fmem_data[7]), .ZN(n1908) );
  OAI22_X1 U1926 ( .A1(n1750), .A2(n1908), .B1(n1909), .B2(n1701), .ZN(n1957)
         );
  XNOR2_X1 U1927 ( .A(n1837), .B(fmem_data[3]), .ZN(n1727) );
  OAI22_X1 U1928 ( .A1(n1702), .A2(n1727), .B1(n1891), .B2(n1703), .ZN(n1956)
         );
  XNOR2_X1 U1929 ( .A(n1728), .B(fmem_data[1]), .ZN(n1729) );
  OAI22_X1 U1930 ( .A1(n1914), .A2(n1729), .B1(n1912), .B2(n1704), .ZN(n1955)
         );
  FA_X1 U1931 ( .A(n1710), .B(n1709), .CI(n1708), .CO(n1676), .S(n1739) );
  NAND2_X1 U1932 ( .A1(n1742), .A2(n1376), .ZN(n1712) );
  NOR2_X1 U1933 ( .A1(n2018), .A2(n2153), .ZN(n2294) );
  XNOR2_X1 U1934 ( .A(n1714), .B(n1713), .ZN(n1716) );
  FA_X1 U1935 ( .A(n1719), .B(n1718), .CI(n1717), .CO(n1689), .S(n1997) );
  XNOR2_X1 U1936 ( .A(n1721), .B(n1720), .ZN(n1722) );
  XNOR2_X1 U1937 ( .A(n1723), .B(n1722), .ZN(n1979) );
  FA_X1 U1938 ( .A(n1726), .B(n1725), .CI(n1724), .CO(n1713), .S(n1978) );
  XNOR2_X1 U1939 ( .A(n1837), .B(fmem_data[2]), .ZN(n1890) );
  OAI22_X1 U1940 ( .A1(n1890), .A2(n1893), .B1(n1891), .B2(n1727), .ZN(n1879)
         );
  XNOR2_X1 U1941 ( .A(\DP_OP_485J1_122_4413/n1204 ), .B(n1728), .ZN(n1730) );
  OAI22_X1 U1942 ( .A1(n1914), .A2(n1730), .B1(n1912), .B2(n1729), .ZN(n1878)
         );
  OR2_X1 U1943 ( .A1(n1879), .A2(n1878), .ZN(n1967) );
  XNOR2_X1 U1944 ( .A(n1745), .B(fmem_data[5]), .ZN(n1884) );
  OAI22_X1 U1945 ( .A1(n1887), .A2(n1884), .B1(n1885), .B2(n1731), .ZN(n1966)
         );
  XNOR2_X1 U1946 ( .A(n1733), .B(n1732), .ZN(n1965) );
  NAND2_X1 U1947 ( .A1(n1735), .A2(n1734), .ZN(n1736) );
  NAND2_X1 U1948 ( .A1(n1998), .A2(n1736), .ZN(n1738) );
  XNOR2_X1 U1949 ( .A(n1740), .B(n1739), .ZN(n1741) );
  XNOR2_X1 U1950 ( .A(n1742), .B(n1741), .ZN(n2020) );
  NOR2_X1 U1951 ( .A1(n2019), .A2(n2020), .ZN(n2368) );
  NOR2_X1 U1952 ( .A1(n2294), .A2(n2368), .ZN(n1743) );
  XNOR2_X1 U1953 ( .A(n1866), .B(fmem_data[1]), .ZN(n1746) );
  XNOR2_X1 U1954 ( .A(n1745), .B(fmem_data[2]), .ZN(n1841) );
  OAI22_X1 U1955 ( .A1(n1887), .A2(n1746), .B1(n1885), .B2(n1841), .ZN(n1836)
         );
  INV_X1 U1956 ( .A(n1891), .ZN(n1744) );
  AND2_X1 U1957 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1744), .ZN(n1835) );
  XNOR2_X1 U1958 ( .A(n1869), .B(fmem_data[5]), .ZN(n1748) );
  XNOR2_X1 U1959 ( .A(n1869), .B(fmem_data[6]), .ZN(n1829) );
  OAI22_X1 U1960 ( .A1(n1779), .A2(n1748), .B1(n1829), .B2(n1882), .ZN(n1834)
         );
  XNOR2_X1 U1961 ( .A(\DP_OP_485J1_122_4413/n1204 ), .B(n1745), .ZN(n1747) );
  OAI22_X1 U1962 ( .A1(n1887), .A2(n1747), .B1(n1885), .B2(n1746), .ZN(n1760)
         );
  NAND2_X2 U1963 ( .A1(xmem_data[1]), .A2(n3328), .ZN(n1906) );
  XNOR2_X1 U1964 ( .A(xmem_data[1]), .B(fmem_data[6]), .ZN(n1770) );
  XNOR2_X1 U1965 ( .A(xmem_data[1]), .B(fmem_data[7]), .ZN(n1752) );
  OAI22_X1 U1966 ( .A1(n1906), .A2(n1770), .B1(n1752), .B2(n3328), .ZN(n1759)
         );
  XNOR2_X1 U1967 ( .A(n1869), .B(fmem_data[4]), .ZN(n1755) );
  OR2_X1 U1968 ( .A1(n1791), .A2(n1799), .ZN(n1880) );
  OAI22_X1 U1969 ( .A1(n1748), .A2(n1882), .B1(n1755), .B2(n1880), .ZN(n1758)
         );
  INV_X1 U1970 ( .A(n1894), .ZN(n1769) );
  XNOR2_X1 U1971 ( .A(n1894), .B(fmem_data[2]), .ZN(n1754) );
  XNOR2_X1 U1972 ( .A(n1894), .B(fmem_data[3]), .ZN(n1751) );
  OAI22_X1 U1973 ( .A1(n1833), .A2(n1754), .B1(n1909), .B2(n1751), .ZN(n1757)
         );
  OR2_X1 U1974 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n3329), .ZN(n1749) );
  OAI22_X1 U1975 ( .A1(n1887), .A2(n3329), .B1(n1749), .B2(n1885), .ZN(n1756)
         );
  XNOR2_X1 U1976 ( .A(n1894), .B(fmem_data[4]), .ZN(n1832) );
  OAI22_X1 U1977 ( .A1(n1911), .A2(n1751), .B1(n1909), .B2(n1832), .ZN(n1846)
         );
  XNOR2_X1 U1978 ( .A(xmem_data[1]), .B(fmem_data[8]), .ZN(n1840) );
  OAI22_X1 U1979 ( .A1(n1906), .A2(n1752), .B1(n1840), .B2(n3328), .ZN(n1845)
         );
  XNOR2_X1 U1980 ( .A(n1846), .B(n1845), .ZN(n1753) );
  XNOR2_X1 U1981 ( .A(n1844), .B(n1753), .ZN(n1850) );
  XNOR2_X1 U1982 ( .A(n1894), .B(fmem_data[1]), .ZN(n1775) );
  OAI22_X1 U1983 ( .A1(n1911), .A2(n1775), .B1(n1909), .B2(n1754), .ZN(n1766)
         );
  AND2_X1 U1984 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1444), .ZN(n1765) );
  XNOR2_X1 U1985 ( .A(n1869), .B(fmem_data[3]), .ZN(n1767) );
  OAI22_X1 U1986 ( .A1(n1767), .A2(n1779), .B1(n1755), .B2(n1882), .ZN(n1764)
         );
  HA_X1 U1987 ( .A(n1757), .B(n1756), .CO(n1844), .S(n1762) );
  FA_X1 U1988 ( .A(n1760), .B(n1759), .CI(n1758), .CO(n1851), .S(n1761) );
  FA_X1 U1989 ( .A(n1763), .B(n1762), .CI(n1761), .CO(n1822), .S(n1825) );
  FA_X1 U1990 ( .A(n1766), .B(n1765), .CI(n1764), .CO(n1763), .S(n1815) );
  XNOR2_X1 U1991 ( .A(n1869), .B(fmem_data[2]), .ZN(n1780) );
  OAI22_X1 U1992 ( .A1(n1767), .A2(n1882), .B1(n1780), .B2(n1880), .ZN(n1778)
         );
  OR2_X1 U1993 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1769), .ZN(n1768) );
  OAI22_X1 U1994 ( .A1(n1833), .A2(n1769), .B1(n1768), .B2(n1909), .ZN(n1777)
         );
  XNOR2_X1 U1995 ( .A(xmem_data[1]), .B(fmem_data[5]), .ZN(n1774) );
  OAI22_X1 U1996 ( .A1(n1906), .A2(n1774), .B1(n1770), .B2(n3328), .ZN(n1812)
         );
  NOR2_X1 U1997 ( .A1(n1825), .A2(n1824), .ZN(n2169) );
  INV_X1 U1998 ( .A(n2169), .ZN(n2356) );
  NAND2_X1 U1999 ( .A1(n2186), .A2(n2356), .ZN(n1828) );
  XNOR2_X1 U2000 ( .A(xmem_data[1]), .B(fmem_data[4]), .ZN(n1784) );
  OAI22_X1 U2001 ( .A1(n1906), .A2(n1784), .B1(n1774), .B2(n3328), .ZN(n1818)
         );
  XNOR2_X1 U2002 ( .A(\DP_OP_485J1_122_4413/n1204 ), .B(n1894), .ZN(n1776) );
  OAI22_X1 U2003 ( .A1(n1911), .A2(n1776), .B1(n1909), .B2(n1775), .ZN(n1817)
         );
  HA_X1 U2004 ( .A(n1778), .B(n1777), .CO(n1813), .S(n1816) );
  XNOR2_X1 U2005 ( .A(n1869), .B(fmem_data[1]), .ZN(n1792) );
  OR2_X1 U2006 ( .A1(n1792), .A2(n1779), .ZN(n1782) );
  OR2_X1 U2007 ( .A1(n1780), .A2(n1882), .ZN(n1781) );
  NAND2_X1 U2008 ( .A1(n1782), .A2(n1781), .ZN(n1790) );
  INV_X1 U2009 ( .A(n1909), .ZN(n1783) );
  AND2_X1 U2010 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1783), .ZN(n1787) );
  XNOR2_X1 U2011 ( .A(xmem_data[1]), .B(fmem_data[3]), .ZN(n1797) );
  OAI22_X1 U2012 ( .A1(n1906), .A2(n1797), .B1(n1784), .B2(n3328), .ZN(n1788)
         );
  NOR2_X1 U2013 ( .A1(n1811), .A2(n1810), .ZN(n2338) );
  XNOR2_X1 U2014 ( .A(\DP_OP_485J1_122_4413/n1204 ), .B(n1869), .ZN(n1793) );
  OR2_X1 U2015 ( .A1(n1791), .A2(n1799), .ZN(n1871) );
  OAI22_X1 U2016 ( .A1(n1793), .A2(n1871), .B1(n1792), .B2(n1882), .ZN(n1796)
         );
  OR2_X1 U2017 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1352), .ZN(n1794) );
  OAI22_X1 U2018 ( .A1(n1794), .A2(n1882), .B1(n1352), .B2(n1871), .ZN(n1795)
         );
  OR2_X1 U2019 ( .A1(n1808), .A2(n1807), .ZN(n2180) );
  HA_X1 U2020 ( .A(n1796), .B(n1795), .CO(n1807), .S(n1806) );
  XNOR2_X1 U2021 ( .A(xmem_data[1]), .B(fmem_data[2]), .ZN(n1798) );
  OAI22_X1 U2022 ( .A1(n1906), .A2(n1798), .B1(n1797), .B2(n3328), .ZN(n1805)
         );
  NOR2_X1 U2023 ( .A1(n1806), .A2(n1805), .ZN(n2331) );
  XNOR2_X1 U2024 ( .A(xmem_data[1]), .B(fmem_data[1]), .ZN(n1801) );
  OAI22_X1 U2025 ( .A1(n1906), .A2(n1801), .B1(n1798), .B2(n3328), .ZN(n1803)
         );
  AND2_X1 U2026 ( .A1(n1799), .A2(\DP_OP_485J1_122_4413/n1204 ), .ZN(n1802) );
  OR2_X1 U2027 ( .A1(n1803), .A2(n1802), .ZN(n2307) );
  OR2_X1 U2028 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n3330), .ZN(n1800) );
  NAND2_X1 U2029 ( .A1(n1800), .A2(n1906), .ZN(n2301) );
  OAI22_X1 U2030 ( .A1(n1906), .A2(\DP_OP_485J1_122_4413/n1204 ), .B1(n1801), 
        .B2(n3328), .ZN(n2300) );
  NAND2_X1 U2031 ( .A1(n2301), .A2(n2300), .ZN(n2302) );
  INV_X1 U2032 ( .A(n2302), .ZN(n2308) );
  NAND2_X1 U2033 ( .A1(n1803), .A2(n1802), .ZN(n2306) );
  INV_X1 U2034 ( .A(n2306), .ZN(n1804) );
  AOI21_X1 U2035 ( .B1(n2307), .B2(n2308), .A(n1804), .ZN(n2334) );
  NAND2_X1 U2036 ( .A1(n1806), .A2(n1805), .ZN(n2332) );
  OAI21_X1 U2037 ( .B1(n2331), .B2(n2334), .A(n2332), .ZN(n2181) );
  INV_X1 U2038 ( .A(n2179), .ZN(n1809) );
  AOI21_X1 U2039 ( .B1(n2180), .B2(n2181), .A(n1809), .ZN(n2342) );
  NAND2_X1 U2040 ( .A1(n1811), .A2(n1810), .ZN(n2339) );
  OAI21_X1 U2041 ( .B1(n2338), .B2(n2342), .A(n2339), .ZN(n2073) );
  FA_X1 U2042 ( .A(n1818), .B(n1817), .CI(n1816), .CO(n1819), .S(n1811) );
  OR2_X1 U2043 ( .A1(n1820), .A2(n1819), .ZN(n2072) );
  NAND2_X1 U2044 ( .A1(n1820), .A2(n1819), .ZN(n2071) );
  INV_X1 U2045 ( .A(n2071), .ZN(n1821) );
  NAND2_X1 U2046 ( .A1(n1823), .A2(n1822), .ZN(n2185) );
  NAND2_X1 U2047 ( .A1(n1825), .A2(n1824), .ZN(n2355) );
  NAND2_X1 U2048 ( .A1(n2185), .A2(n2355), .ZN(n1826) );
  NAND2_X1 U2049 ( .A1(n2186), .A2(n1826), .ZN(n1827) );
  OAI21_X1 U2050 ( .B1(n1828), .B2(n2358), .A(n1827), .ZN(n1858) );
  XNOR2_X1 U2051 ( .A(n1869), .B(fmem_data[7]), .ZN(n1870) );
  OAI22_X1 U2052 ( .A1(n1829), .A2(n1871), .B1(n1870), .B2(n1882), .ZN(n1860)
         );
  XNOR2_X1 U2053 ( .A(\DP_OP_485J1_122_4413/n1204 ), .B(n1837), .ZN(n1830) );
  XNOR2_X1 U2054 ( .A(n1837), .B(fmem_data[1]), .ZN(n1892) );
  OAI22_X1 U2055 ( .A1(n1831), .A2(n1830), .B1(n1891), .B2(n1892), .ZN(n1859)
         );
  XNOR2_X1 U2056 ( .A(n1894), .B(fmem_data[5]), .ZN(n1895) );
  OAI22_X1 U2057 ( .A1(n1833), .A2(n1832), .B1(n1909), .B2(n1895), .ZN(n1917)
         );
  FA_X1 U2058 ( .A(n1836), .B(n1835), .CI(n1834), .CO(n1916), .S(n1852) );
  INV_X1 U2059 ( .A(n1837), .ZN(n1839) );
  OR2_X1 U2060 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n1839), .ZN(n1838) );
  OAI22_X1 U2061 ( .A1(n1893), .A2(n1839), .B1(n1838), .B2(n1891), .ZN(n1862)
         );
  XNOR2_X1 U2062 ( .A(xmem_data[1]), .B(fmem_data[9]), .ZN(n1896) );
  OAI22_X1 U2063 ( .A1(n1906), .A2(n1840), .B1(n1896), .B2(n3328), .ZN(n1861)
         );
  XNOR2_X1 U2064 ( .A(n1866), .B(fmem_data[3]), .ZN(n1867) );
  OAI22_X1 U2065 ( .A1(n1887), .A2(n1841), .B1(n1885), .B2(n1867), .ZN(n1863)
         );
  XNOR2_X1 U2066 ( .A(n1842), .B(n1863), .ZN(n1930) );
  INV_X1 U2067 ( .A(n1856), .ZN(n1854) );
  FA_X1 U2068 ( .A(n1852), .B(n1851), .CI(n1850), .CO(n1855), .S(n1823) );
  INV_X1 U2069 ( .A(n1855), .ZN(n1853) );
  NAND2_X1 U2070 ( .A1(n1854), .A2(n1853), .ZN(n2362) );
  NAND2_X1 U2071 ( .A1(n1856), .A2(n1855), .ZN(n2361) );
  INV_X1 U2072 ( .A(n2361), .ZN(n1857) );
  AOI21_X1 U2073 ( .B1(n1858), .B2(n2362), .A(n1857), .ZN(n2148) );
  HA_X1 U2074 ( .A(n1860), .B(n1859), .CO(n1922), .S(n1918) );
  OAI21_X1 U2075 ( .B1(n1862), .B2(n1863), .A(n1861), .ZN(n1865) );
  NAND2_X1 U2076 ( .A1(n1863), .A2(n1862), .ZN(n1864) );
  NAND2_X1 U2077 ( .A1(n1865), .A2(n1864), .ZN(n1923) );
  OR2_X1 U2078 ( .A1(n1922), .A2(n1923), .ZN(n1875) );
  XNOR2_X1 U2079 ( .A(n1866), .B(fmem_data[4]), .ZN(n1886) );
  OAI22_X1 U2080 ( .A1(n1887), .A2(n1867), .B1(n1885), .B2(n1886), .ZN(n1902)
         );
  NAND2_X1 U2081 ( .A1(n1868), .A2(\DP_OP_485J1_122_4413/n1204 ), .ZN(n1897)
         );
  INV_X1 U2082 ( .A(n1897), .ZN(n1901) );
  XNOR2_X1 U2083 ( .A(n1902), .B(n1901), .ZN(n1874) );
  XNOR2_X1 U2084 ( .A(n1869), .B(fmem_data[8]), .ZN(n1881) );
  OR2_X1 U2085 ( .A1(n1881), .A2(n1882), .ZN(n1873) );
  NAND2_X1 U2086 ( .A1(n1873), .A2(n1872), .ZN(n1900) );
  XNOR2_X1 U2087 ( .A(n1874), .B(n1900), .ZN(n1925) );
  NAND2_X1 U2088 ( .A1(n1875), .A2(n1925), .ZN(n1877) );
  NAND2_X1 U2089 ( .A1(n1877), .A2(n1876), .ZN(n1974) );
  OR2_X1 U2090 ( .A1(n1881), .A2(n1880), .ZN(n1945) );
  OR2_X1 U2091 ( .A1(n1883), .A2(n1882), .ZN(n1946) );
  NAND2_X1 U2092 ( .A1(n1945), .A2(n1946), .ZN(n1888) );
  OAI22_X1 U2093 ( .A1(n1887), .A2(n1886), .B1(n1885), .B2(n1884), .ZN(n1948)
         );
  XNOR2_X1 U2094 ( .A(n1888), .B(n1948), .ZN(n1889) );
  XNOR2_X1 U2095 ( .A(n1952), .B(n1889), .ZN(n1973) );
  XNOR2_X1 U2096 ( .A(n1974), .B(n1973), .ZN(n1915) );
  OAI22_X1 U2097 ( .A1(n1893), .A2(n1892), .B1(n1891), .B2(n1890), .ZN(n1921)
         );
  XNOR2_X1 U2098 ( .A(n1894), .B(fmem_data[6]), .ZN(n1910) );
  OAI22_X1 U2099 ( .A1(n1911), .A2(n1895), .B1(n1909), .B2(n1910), .ZN(n1920)
         );
  XNOR2_X1 U2100 ( .A(xmem_data[1]), .B(fmem_data[19]), .ZN(n1905) );
  OAI22_X1 U2101 ( .A1(n1906), .A2(n1896), .B1(n1905), .B2(n3328), .ZN(n1919)
         );
  INV_X1 U2102 ( .A(n1902), .ZN(n1898) );
  NAND2_X1 U2103 ( .A1(n1898), .A2(n1897), .ZN(n1899) );
  NAND2_X1 U2104 ( .A1(n1900), .A2(n1899), .ZN(n1904) );
  NAND2_X1 U2105 ( .A1(n1902), .A2(n1901), .ZN(n1903) );
  NAND2_X1 U2106 ( .A1(n1904), .A2(n1903), .ZN(n1963) );
  AOI21_X1 U2107 ( .B1(n1906), .B2(n3328), .A(n1905), .ZN(n1907) );
  INV_X1 U2108 ( .A(n1907), .ZN(n1960) );
  OAI22_X1 U2109 ( .A1(n1911), .A2(n1910), .B1(n1909), .B2(n1908), .ZN(n1959)
         );
  OR2_X1 U2110 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(n3391), .ZN(n1913) );
  OAI22_X1 U2111 ( .A1(n1914), .A2(n3391), .B1(n1913), .B2(n1912), .ZN(n1958)
         );
  XNOR2_X1 U2112 ( .A(n1915), .B(n1971), .ZN(n1943) );
  FA_X1 U2113 ( .A(n1918), .B(n1917), .CI(n1916), .CO(n1935), .S(n1929) );
  FA_X1 U2114 ( .A(n1921), .B(n1920), .CI(n1919), .CO(n1964), .S(n1934) );
  XNOR2_X1 U2115 ( .A(n1923), .B(n1922), .ZN(n1924) );
  XNOR2_X1 U2116 ( .A(n1925), .B(n1924), .ZN(n1936) );
  OAI21_X1 U2117 ( .B1(n1935), .B2(n1934), .A(n1936), .ZN(n1927) );
  NAND2_X1 U2118 ( .A1(n1935), .A2(n1934), .ZN(n1926) );
  NAND2_X1 U2119 ( .A1(n1927), .A2(n1926), .ZN(n1942) );
  NOR2_X1 U2120 ( .A1(n1943), .A2(n1942), .ZN(n2168) );
  INV_X1 U2121 ( .A(n2168), .ZN(n2350) );
  INV_X1 U2122 ( .A(n1941), .ZN(n1939) );
  XNOR2_X1 U2123 ( .A(n1935), .B(n1934), .ZN(n1937) );
  XNOR2_X1 U2124 ( .A(n1937), .B(n1936), .ZN(n1940) );
  INV_X1 U2125 ( .A(n1940), .ZN(n1938) );
  NAND2_X1 U2126 ( .A1(n1939), .A2(n1938), .ZN(n2348) );
  NAND2_X1 U2127 ( .A1(n2350), .A2(n2348), .ZN(n2149) );
  NAND2_X1 U2128 ( .A1(n1941), .A2(n1940), .ZN(n2346) );
  NAND2_X1 U2129 ( .A1(n1943), .A2(n1942), .ZN(n2349) );
  OAI21_X1 U2130 ( .B1(n2168), .B2(n2346), .A(n2349), .ZN(n1944) );
  INV_X1 U2131 ( .A(n1944), .ZN(n2172) );
  OAI21_X1 U2132 ( .B1(n2148), .B2(n2149), .A(n2172), .ZN(n2017) );
  AND2_X1 U2133 ( .A1(n1946), .A2(n1945), .ZN(n1949) );
  INV_X1 U2134 ( .A(n1949), .ZN(n1947) );
  NAND2_X1 U2135 ( .A1(n1950), .A2(n1949), .ZN(n1951) );
  NAND2_X1 U2136 ( .A1(n1952), .A2(n1951), .ZN(n1953) );
  NAND2_X1 U2137 ( .A1(n1954), .A2(n1953), .ZN(n1980) );
  FA_X1 U2138 ( .A(n1957), .B(n1956), .CI(n1955), .CO(n1986), .S(n1983) );
  FA_X1 U2139 ( .A(n1960), .B(n1959), .CI(n1958), .CO(n1982), .S(n1962) );
  XNOR2_X1 U2140 ( .A(n1983), .B(n1982), .ZN(n1961) );
  FA_X1 U2141 ( .A(n1964), .B(n1963), .CI(n1962), .CO(n1993), .S(n1971) );
  FA_X1 U2142 ( .A(n1967), .B(n1966), .CI(n1965), .CO(n1977), .S(n1992) );
  XNOR2_X1 U2143 ( .A(n1993), .B(n1992), .ZN(n1968) );
  XNOR2_X1 U2144 ( .A(n1990), .B(n1968), .ZN(n2007) );
  INV_X1 U2145 ( .A(n1974), .ZN(n1970) );
  NAND2_X1 U2146 ( .A1(n1970), .A2(n1969), .ZN(n1972) );
  NAND2_X1 U2147 ( .A1(n1972), .A2(n1971), .ZN(n1976) );
  NAND2_X1 U2148 ( .A1(n1974), .A2(n1973), .ZN(n1975) );
  NAND2_X1 U2149 ( .A1(n1976), .A2(n1975), .ZN(n2006) );
  NOR2_X1 U2150 ( .A1(n2007), .A2(n2006), .ZN(n2175) );
  FA_X1 U2151 ( .A(n1979), .B(n1978), .CI(n1977), .CO(n1996), .S(n2000) );
  OR2_X1 U2152 ( .A1(n1983), .A2(n1982), .ZN(n1981) );
  NAND2_X1 U2153 ( .A1(n1981), .A2(n1980), .ZN(n1985) );
  NAND2_X1 U2154 ( .A1(n1983), .A2(n1982), .ZN(n1984) );
  NAND2_X1 U2155 ( .A1(n1985), .A2(n1984), .ZN(n2002) );
  FA_X1 U2156 ( .A(n1988), .B(n1987), .CI(n1986), .CO(n1715), .S(n2001) );
  XNOR2_X1 U2157 ( .A(n2002), .B(n2001), .ZN(n1989) );
  XNOR2_X1 U2158 ( .A(n2000), .B(n1989), .ZN(n2009) );
  OR2_X1 U2159 ( .A1(n1993), .A2(n1992), .ZN(n1991) );
  NAND2_X1 U2160 ( .A1(n1991), .A2(n1990), .ZN(n1995) );
  NAND2_X1 U2161 ( .A1(n1993), .A2(n1992), .ZN(n1994) );
  NAND2_X1 U2162 ( .A1(n1995), .A2(n1994), .ZN(n2008) );
  OR2_X2 U2163 ( .A1(n2009), .A2(n2008), .ZN(n2314) );
  NAND2_X1 U2164 ( .A1(n1340), .A2(n2314), .ZN(n2005) );
  XNOR2_X1 U2165 ( .A(n1997), .B(n1996), .ZN(n1999) );
  XNOR2_X1 U2166 ( .A(n1999), .B(n1998), .ZN(n2012) );
  NAND2_X1 U2167 ( .A1(n2000), .A2(n1377), .ZN(n2004) );
  NAND2_X1 U2168 ( .A1(n2002), .A2(n2001), .ZN(n2003) );
  NOR2_X1 U2169 ( .A1(n2012), .A2(n2011), .ZN(n2324) );
  NOR2_X1 U2170 ( .A1(n2005), .A2(n2324), .ZN(n2016) );
  NAND2_X1 U2171 ( .A1(n2007), .A2(n2006), .ZN(n2150) );
  INV_X1 U2172 ( .A(n2150), .ZN(n2010) );
  AND2_X1 U2173 ( .A1(n2009), .A2(n2008), .ZN(n2151) );
  AOI21_X1 U2174 ( .B1(n2314), .B2(n2010), .A(n2151), .ZN(n2014) );
  NOR2_X1 U2175 ( .A1(n2012), .A2(n2011), .ZN(n2013) );
  NAND2_X1 U2176 ( .A1(n2012), .A2(n2011), .ZN(n2325) );
  OAI21_X1 U2177 ( .B1(n2014), .B2(n2013), .A(n2325), .ZN(n2015) );
  AOI21_X1 U2178 ( .B1(n2017), .B2(n2016), .A(n2015), .ZN(n2367) );
  NOR2_X1 U2179 ( .A1(n2018), .A2(n2153), .ZN(n2025) );
  NAND2_X1 U2180 ( .A1(n2020), .A2(n2019), .ZN(n2369) );
  FA_X1 U2181 ( .A(n1342), .B(n2022), .CI(n2021), .CO(n2026), .S(n2154) );
  NAND2_X1 U2182 ( .A1(n2154), .A2(n2153), .ZN(n2024) );
  OAI21_X1 U2183 ( .B1(n2025), .B2(n2369), .A(n2024), .ZN(n2032) );
  NAND2_X1 U2184 ( .A1(n2027), .A2(n2026), .ZN(n2384) );
  NAND2_X1 U2185 ( .A1(n2029), .A2(n2028), .ZN(n2393) );
  OAI21_X1 U2186 ( .B1(n2392), .B2(n2384), .A(n2393), .ZN(n2030) );
  AOI21_X1 U2187 ( .B1(n2031), .B2(n2032), .A(n2030), .ZN(n2033) );
  OAI21_X1 U2188 ( .B1(n2034), .B2(n2367), .A(n2033), .ZN(n2792) );
  NAND2_X1 U2189 ( .A1(n2788), .A2(n2786), .ZN(n2079) );
  NAND2_X1 U2190 ( .A1(n2035), .A2(n2080), .ZN(n2036) );
  OAI21_X1 U2191 ( .B1(n2037), .B2(n2079), .A(n2036), .ZN(n2046) );
  NAND2_X1 U2192 ( .A1(n2039), .A2(n2038), .ZN(n2044) );
  INV_X1 U2193 ( .A(n1343), .ZN(n2043) );
  NAND2_X1 U2194 ( .A1(n2041), .A2(n1343), .ZN(n2042) );
  OAI21_X1 U2195 ( .B1(n2044), .B2(n2043), .A(n2042), .ZN(n2045) );
  AOI21_X1 U2196 ( .B1(n2047), .B2(n2046), .A(n2045), .ZN(n2066) );
  NAND2_X1 U2197 ( .A1(n2049), .A2(n2048), .ZN(n2061) );
  AND2_X1 U2198 ( .A1(n2051), .A2(n2050), .ZN(n2053) );
  NAND2_X1 U2199 ( .A1(n2053), .A2(n2052), .ZN(n2059) );
  HA_X1 U2200 ( .A(n2097), .B(n2098), .CO(n2055), .S(n2050) );
  NAND2_X1 U2201 ( .A1(n2055), .A2(n2054), .ZN(n2058) );
  INV_X1 U2202 ( .A(n2056), .ZN(n2057) );
  OAI211_X1 U2203 ( .C1(n2061), .C2(n2060), .A(n2059), .B(n1386), .ZN(n2062)
         );
  NAND2_X1 U2204 ( .A1(n2063), .A2(n2062), .ZN(n2064) );
  OAI21_X1 U2205 ( .B1(n2066), .B2(n2065), .A(n2064), .ZN(n2067) );
  AOI21_X1 U2206 ( .B1(n2068), .B2(n2792), .A(n2067), .ZN(n2793) );
  NAND2_X1 U2207 ( .A1(m_valid_y), .A2(m_ready_y), .ZN(n2820) );
  INV_X1 U2208 ( .A(reset), .ZN(n2815) );
  NAND2_X1 U2209 ( .A1(n2820), .A2(n2815), .ZN(n3307) );
  INV_X1 U2210 ( .A(n3307), .ZN(n2070) );
  NAND2_X1 U2211 ( .A1(n3367), .A2(conv_pre_start), .ZN(n2818) );
  NOR2_X1 U2212 ( .A1(n2818), .A2(n3368), .ZN(n2069) );
  NAND2_X1 U2213 ( .A1(n2070), .A2(n2069), .ZN(n2164) );
  NOR2_X1 U2214 ( .A1(n2793), .A2(n2164), .ZN(n2287) );
  BUF_X2 U2215 ( .A(n2287), .Z(n2397) );
  NAND2_X1 U2216 ( .A1(n2072), .A2(n2071), .ZN(n2074) );
  XNOR2_X1 U2217 ( .A(n2074), .B(n1341), .ZN(n2075) );
  NAND2_X1 U2218 ( .A1(n2397), .A2(n2075), .ZN(n2166) );
  XNOR2_X1 U2219 ( .A(n2076), .B(n2089), .ZN(n2083) );
  NAND2_X1 U2220 ( .A1(n2077), .A2(n2786), .ZN(n2082) );
  NOR2_X1 U2221 ( .A1(n2083), .A2(n2082), .ZN(n2086) );
  XNOR2_X1 U2222 ( .A(n2077), .B(n2786), .ZN(n2081) );
  NOR2_X1 U2223 ( .A1(n2081), .A2(n2080), .ZN(n2078) );
  NOR2_X1 U2224 ( .A1(n2086), .A2(n2078), .ZN(n2145) );
  OAI21_X1 U2225 ( .B1(n2143), .B2(n2393), .A(n2079), .ZN(n2088) );
  NAND2_X1 U2226 ( .A1(n2081), .A2(n2080), .ZN(n2085) );
  NAND2_X1 U2227 ( .A1(n2083), .A2(n2082), .ZN(n2084) );
  OAI21_X1 U2228 ( .B1(n2086), .B2(n2085), .A(n2084), .ZN(n2087) );
  AOI21_X1 U2229 ( .B1(n2145), .B2(n2088), .A(n2087), .ZN(n2141) );
  OR2_X1 U2230 ( .A1(n2090), .A2(n2089), .ZN(n2105) );
  XNOR2_X1 U2231 ( .A(n2092), .B(n2093), .ZN(n2104) );
  NOR2_X1 U2232 ( .A1(n2105), .A2(n2104), .ZN(n2094) );
  XNOR2_X1 U2233 ( .A(n2091), .B(n2095), .ZN(n2107) );
  OR2_X1 U2234 ( .A1(n2093), .A2(n2092), .ZN(n2106) );
  NOR2_X1 U2235 ( .A1(n2107), .A2(n2106), .ZN(n2109) );
  NOR2_X1 U2236 ( .A1(n2094), .A2(n2109), .ZN(n2103) );
  OR2_X1 U2237 ( .A1(n2096), .A2(n2095), .ZN(n2112) );
  XNOR2_X1 U2238 ( .A(n2098), .B(n2097), .ZN(n2111) );
  OR2_X1 U2239 ( .A1(n2112), .A2(n2111), .ZN(n2099) );
  OR2_X1 U2240 ( .A1(n2098), .A2(n2097), .ZN(n2116) );
  NAND2_X1 U2241 ( .A1(n2099), .A2(n2116), .ZN(n2102) );
  OR2_X1 U2242 ( .A1(n2119), .A2(n2118), .ZN(n2100) );
  OR2_X1 U2243 ( .A1(n2121), .A2(n2120), .ZN(n2124) );
  NAND2_X1 U2244 ( .A1(n2100), .A2(n2124), .ZN(n2127) );
  NOR2_X1 U2245 ( .A1(n1356), .A2(n2127), .ZN(n2101) );
  NOR2_X1 U2246 ( .A1(n2129), .A2(n2128), .ZN(n2130) );
  NOR2_X1 U2247 ( .A1(n1355), .A2(n2130), .ZN(n2132) );
  NAND2_X1 U2248 ( .A1(n2101), .A2(n2132), .ZN(n2135) );
  NOR2_X1 U2249 ( .A1(n2102), .A2(n2135), .ZN(n2139) );
  NAND2_X1 U2250 ( .A1(n2103), .A2(n2139), .ZN(n2146) );
  NAND2_X1 U2251 ( .A1(n2105), .A2(n2104), .ZN(n2110) );
  NAND2_X1 U2252 ( .A1(n2107), .A2(n2106), .ZN(n2108) );
  OAI21_X1 U2253 ( .B1(n2110), .B2(n2109), .A(n2108), .ZN(n2138) );
  AND2_X1 U2254 ( .A1(n2112), .A2(n2111), .ZN(n2117) );
  XNOR2_X1 U2255 ( .A(n2114), .B(n2113), .ZN(n2115) );
  AOI21_X1 U2256 ( .B1(n2117), .B2(n2116), .A(n2115), .ZN(n2136) );
  XNOR2_X1 U2257 ( .A(n2121), .B(n2120), .ZN(n2125) );
  AOI21_X1 U2258 ( .B1(n2125), .B2(n2124), .A(n1385), .ZN(n2126) );
  OAI21_X1 U2259 ( .B1(n2127), .B2(n1354), .A(n2126), .ZN(n2133) );
  NOR2_X1 U2260 ( .A1(n1353), .A2(n2130), .ZN(n2131) );
  AOI21_X1 U2261 ( .B1(n2133), .B2(n2132), .A(n2131), .ZN(n2134) );
  OAI21_X1 U2262 ( .B1(n2136), .B2(n2135), .A(n2134), .ZN(n2137) );
  AOI21_X1 U2263 ( .B1(n2139), .B2(n2138), .A(n2137), .ZN(n2140) );
  OAI21_X1 U2264 ( .B1(n2141), .B2(n2146), .A(n2140), .ZN(n2142) );
  INV_X1 U2265 ( .A(n2142), .ZN(n2163) );
  NOR2_X1 U2266 ( .A1(n2392), .A2(n2143), .ZN(n2144) );
  NAND2_X1 U2267 ( .A1(n2145), .A2(n2144), .ZN(n2147) );
  NOR2_X1 U2268 ( .A1(n2147), .A2(n2146), .ZN(n2161) );
  OAI21_X1 U2269 ( .B1(n2148), .B2(n2149), .A(n2172), .ZN(n2289) );
  INV_X1 U2270 ( .A(n2314), .ZN(n2152) );
  NOR2_X1 U2271 ( .A1(n2175), .A2(n2152), .ZN(n2319) );
  INV_X1 U2272 ( .A(n2151), .ZN(n2313) );
  OAI21_X1 U2273 ( .B1(n2152), .B2(n2312), .A(n2313), .ZN(n2320) );
  AOI21_X1 U2274 ( .B1(n2289), .B2(n2319), .A(n2320), .ZN(n2159) );
  NOR2_X1 U2275 ( .A1(n2324), .A2(n2368), .ZN(n2291) );
  NOR2_X1 U2276 ( .A1(n2294), .A2(n1344), .ZN(n2156) );
  NAND2_X1 U2277 ( .A1(n2291), .A2(n2156), .ZN(n2158) );
  OAI21_X1 U2278 ( .B1(n2368), .B2(n2325), .A(n2369), .ZN(n2290) );
  NAND2_X1 U2279 ( .A1(n2154), .A2(n2153), .ZN(n2375) );
  OAI21_X1 U2280 ( .B1(n1344), .B2(n2375), .A(n2384), .ZN(n2155) );
  AOI21_X1 U2281 ( .B1(n2290), .B2(n2156), .A(n2155), .ZN(n2157) );
  OAI21_X1 U2282 ( .B1(n2159), .B2(n2158), .A(n2157), .ZN(n2160) );
  NAND2_X1 U2283 ( .A1(n2161), .A2(n2160), .ZN(n2162) );
  NAND2_X1 U2284 ( .A1(n2163), .A2(n2162), .ZN(n2794) );
  INV_X1 U2285 ( .A(n2164), .ZN(n2796) );
  NAND2_X2 U2286 ( .A1(n2794), .A2(n2796), .ZN(n2399) );
  NAND2_X1 U2287 ( .A1(n2818), .A2(\ctrl_conv_output_inst/conv_start_accum ), 
        .ZN(n2165) );
  NAND3_X1 U2288 ( .A1(n2166), .A2(n2399), .A3(n1357), .ZN(n904) );
  NOR2_X1 U2289 ( .A1(n2168), .A2(n2167), .ZN(n2174) );
  OAI21_X1 U2290 ( .B1(n2358), .B2(n2169), .A(n2355), .ZN(n2188) );
  AOI21_X1 U2291 ( .B1(n2188), .B2(n2186), .A(n2170), .ZN(n2364) );
  INV_X1 U2292 ( .A(n2362), .ZN(n2171) );
  OAI21_X1 U2293 ( .B1(n2364), .B2(n2171), .A(n2361), .ZN(n2191) );
  AOI21_X1 U2294 ( .B1(n2174), .B2(n2191), .A(n2173), .ZN(n2323) );
  NAND2_X1 U2295 ( .A1(n1340), .A2(n2312), .ZN(n2176) );
  XOR2_X1 U2296 ( .A(n2323), .B(n2176), .Z(n2177) );
  NAND2_X1 U2297 ( .A1(n2397), .A2(n2177), .ZN(n2178) );
  NAND3_X1 U2298 ( .A1(n2178), .A2(n2399), .A3(n1358), .ZN(n898) );
  NAND2_X1 U2299 ( .A1(n2180), .A2(n2179), .ZN(n2182) );
  XNOR2_X1 U2300 ( .A(n2182), .B(n2181), .ZN(n2183) );
  NAND2_X1 U2301 ( .A1(n2397), .A2(n2183), .ZN(n2184) );
  NAND3_X1 U2302 ( .A1(n2184), .A2(n2399), .A3(n1359), .ZN(n906) );
  NAND2_X1 U2303 ( .A1(n2186), .A2(n2185), .ZN(n2187) );
  XNOR2_X1 U2304 ( .A(n2188), .B(n2187), .ZN(n2189) );
  NAND2_X1 U2305 ( .A1(n2397), .A2(n2189), .ZN(n2190) );
  NAND3_X1 U2306 ( .A1(n2190), .A2(n2399), .A3(n1360), .ZN(n902) );
  INV_X1 U2307 ( .A(n2191), .ZN(n2345) );
  NAND2_X1 U2308 ( .A1(n2348), .A2(n2346), .ZN(n2192) );
  XOR2_X1 U2309 ( .A(n2345), .B(n2192), .Z(n2193) );
  NAND2_X1 U2310 ( .A1(n2397), .A2(n2193), .ZN(n2194) );
  NAND3_X1 U2311 ( .A1(n2194), .A2(n2399), .A3(n1361), .ZN(n900) );
  NAND2_X1 U2312 ( .A1(xmem_addr[0]), .A2(xmem_addr[1]), .ZN(n3184) );
  OR2_X1 U2313 ( .A1(n3340), .A2(n3184), .ZN(n2830) );
  NOR2_X2 U2314 ( .A1(n3335), .A2(n2830), .ZN(n2835) );
  NAND2_X1 U2315 ( .A1(xmem_addr[0]), .A2(n3345), .ZN(n3137) );
  AOI22_X1 U2316 ( .A1(n2835), .A2(\xmem_inst/mem[15][19] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][19] ), .ZN(n2199) );
  NOR3_X1 U2317 ( .A1(n3184), .A2(n3340), .A3(xmem_addr[3]), .ZN(n2831) );
  NAND2_X1 U2318 ( .A1(xmem_addr[1]), .A2(n3338), .ZN(n3160) );
  NOR2_X2 U2319 ( .A1(n3334), .A2(n3160), .ZN(n3253) );
  AOI22_X1 U2320 ( .A1(n2575), .A2(\xmem_inst/mem[7][19] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][19] ), .ZN(n2198) );
  NOR2_X1 U2321 ( .A1(xmem_addr[2]), .A2(xmem_addr[3]), .ZN(n2817) );
  NAND2_X1 U2322 ( .A1(n2817), .A2(n3334), .ZN(n2195) );
  AOI22_X1 U2323 ( .A1(n2442), .A2(\xmem_inst/mem[3][19] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][19] ), .ZN(n2197) );
  NOR2_X2 U2324 ( .A1(n3160), .A2(n2195), .ZN(n2885) );
  NAND2_X1 U2325 ( .A1(n3338), .A2(n3345), .ZN(n3114) );
  AOI22_X1 U2326 ( .A1(n2885), .A2(\xmem_inst/mem[2][19] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][19] ), .ZN(n2196) );
  NAND4_X1 U2327 ( .A1(n2199), .A2(n2198), .A3(n2197), .A4(n2196), .ZN(n2221)
         );
  NOR2_X1 U2328 ( .A1(n3335), .A2(xmem_addr[2]), .ZN(n3022) );
  INV_X1 U2329 ( .A(n3022), .ZN(n2213) );
  NOR2_X1 U2330 ( .A1(n3340), .A2(xmem_addr[3]), .ZN(n2932) );
  INV_X1 U2331 ( .A(n2932), .ZN(n2206) );
  AOI22_X1 U2332 ( .A1(n2200), .A2(\xmem_inst/mem[8][19] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][19] ), .ZN(n2211) );
  NOR2_X1 U2333 ( .A1(n3340), .A2(n3335), .ZN(n3113) );
  INV_X1 U2334 ( .A(n3113), .ZN(n2215) );
  AOI22_X1 U2335 ( .A1(n2202), .A2(\xmem_inst/mem[14][19] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][19] ), .ZN(n2210) );
  AOI22_X1 U2336 ( .A1(n2447), .A2(\xmem_inst/mem[19][19] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][19] ), .ZN(n2209) );
  AOI22_X1 U2337 ( .A1(n2205), .A2(\xmem_inst/mem[6][19] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][19] ), .ZN(n2208) );
  NAND4_X1 U2338 ( .A1(n2211), .A2(n2210), .A3(n2209), .A4(n2208), .ZN(n2220)
         );
  NOR2_X2 U2339 ( .A1(n3334), .A2(n3114), .ZN(n3207) );
  AOI22_X1 U2340 ( .A1(n3207), .A2(\xmem_inst/mem[16][19] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][19] ), .ZN(n2218) );
  AOI22_X1 U2341 ( .A1(n2214), .A2(\xmem_inst/mem[10][19] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][19] ), .ZN(n2217) );
  NAND2_X1 U2342 ( .A1(n2218), .A2(n2217), .ZN(n2219) );
  AOI22_X1 U2343 ( .A1(n2835), .A2(\xmem_inst/mem[15][17] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][17] ), .ZN(n2225) );
  AOI22_X1 U2344 ( .A1(n2575), .A2(\xmem_inst/mem[7][17] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][17] ), .ZN(n2224) );
  AOI22_X1 U2345 ( .A1(n2442), .A2(\xmem_inst/mem[3][17] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][17] ), .ZN(n2223) );
  AOI22_X1 U2346 ( .A1(n2885), .A2(\xmem_inst/mem[2][17] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][17] ), .ZN(n2222) );
  NAND4_X1 U2347 ( .A1(n2225), .A2(n2224), .A3(n2223), .A4(n2222), .ZN(n2234)
         );
  AOI22_X1 U2348 ( .A1(n2200), .A2(\xmem_inst/mem[8][17] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][17] ), .ZN(n2229) );
  AOI22_X1 U2349 ( .A1(n2202), .A2(\xmem_inst/mem[14][17] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][17] ), .ZN(n2228) );
  AOI22_X1 U2350 ( .A1(n2447), .A2(\xmem_inst/mem[19][17] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][17] ), .ZN(n2227) );
  AOI22_X1 U2351 ( .A1(n2205), .A2(\xmem_inst/mem[6][17] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][17] ), .ZN(n2226) );
  NAND4_X1 U2352 ( .A1(n2229), .A2(n2228), .A3(n2227), .A4(n2226), .ZN(n2233)
         );
  AOI22_X1 U2353 ( .A1(n3207), .A2(\xmem_inst/mem[16][17] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][17] ), .ZN(n2231) );
  AOI22_X1 U2354 ( .A1(n2214), .A2(\xmem_inst/mem[10][17] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][17] ), .ZN(n2230) );
  NAND2_X1 U2355 ( .A1(n2231), .A2(n2230), .ZN(n2232) );
  AOI22_X1 U2356 ( .A1(n2835), .A2(\xmem_inst/mem[15][13] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][13] ), .ZN(n2238) );
  AOI22_X1 U2357 ( .A1(n2575), .A2(\xmem_inst/mem[7][13] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][13] ), .ZN(n2237) );
  AOI22_X1 U2358 ( .A1(n2442), .A2(\xmem_inst/mem[3][13] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][13] ), .ZN(n2236) );
  AOI22_X1 U2359 ( .A1(n2885), .A2(\xmem_inst/mem[2][13] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][13] ), .ZN(n2235) );
  NAND4_X1 U2360 ( .A1(n2238), .A2(n2237), .A3(n2236), .A4(n2235), .ZN(n2247)
         );
  AOI22_X1 U2361 ( .A1(n2200), .A2(\xmem_inst/mem[8][13] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][13] ), .ZN(n2242) );
  AOI22_X1 U2362 ( .A1(n2202), .A2(\xmem_inst/mem[14][13] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][13] ), .ZN(n2241) );
  AOI22_X1 U2363 ( .A1(n2447), .A2(\xmem_inst/mem[19][13] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][13] ), .ZN(n2240) );
  AOI22_X1 U2364 ( .A1(n2205), .A2(\xmem_inst/mem[6][13] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][13] ), .ZN(n2239) );
  NAND4_X1 U2365 ( .A1(n2242), .A2(n2241), .A3(n2240), .A4(n2239), .ZN(n2246)
         );
  AOI22_X1 U2366 ( .A1(n3207), .A2(\xmem_inst/mem[16][13] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][13] ), .ZN(n2244) );
  AOI22_X1 U2367 ( .A1(n2214), .A2(\xmem_inst/mem[10][13] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][13] ), .ZN(n2243) );
  NAND2_X1 U2368 ( .A1(n2244), .A2(n2243), .ZN(n2245) );
  AOI22_X1 U2369 ( .A1(n2835), .A2(\xmem_inst/mem[15][5] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][5] ), .ZN(n2251) );
  AOI22_X1 U2370 ( .A1(n2575), .A2(\xmem_inst/mem[7][5] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][5] ), .ZN(n2250) );
  AOI22_X1 U2371 ( .A1(n2442), .A2(\xmem_inst/mem[3][5] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][5] ), .ZN(n2249) );
  AOI22_X1 U2372 ( .A1(n2885), .A2(\xmem_inst/mem[2][5] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][5] ), .ZN(n2248) );
  NAND4_X1 U2373 ( .A1(n2251), .A2(n2250), .A3(n2249), .A4(n2248), .ZN(n2260)
         );
  AOI22_X1 U2374 ( .A1(n2200), .A2(\xmem_inst/mem[8][5] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][5] ), .ZN(n2255) );
  AOI22_X1 U2375 ( .A1(n2202), .A2(\xmem_inst/mem[14][5] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][5] ), .ZN(n2254) );
  AOI22_X1 U2376 ( .A1(n2447), .A2(\xmem_inst/mem[19][5] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][5] ), .ZN(n2253) );
  AOI22_X1 U2377 ( .A1(n2205), .A2(\xmem_inst/mem[6][5] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][5] ), .ZN(n2252) );
  NAND4_X1 U2378 ( .A1(n2255), .A2(n2254), .A3(n2253), .A4(n2252), .ZN(n2259)
         );
  AOI22_X1 U2379 ( .A1(n3207), .A2(\xmem_inst/mem[16][5] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][5] ), .ZN(n2257) );
  AOI22_X1 U2380 ( .A1(n2214), .A2(\xmem_inst/mem[10][5] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][5] ), .ZN(n2256) );
  NAND2_X1 U2381 ( .A1(n2257), .A2(n2256), .ZN(n2258) );
  AOI22_X1 U2382 ( .A1(n2835), .A2(\xmem_inst/mem[15][7] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][7] ), .ZN(n2264) );
  AOI22_X1 U2383 ( .A1(n2575), .A2(\xmem_inst/mem[7][7] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][7] ), .ZN(n2263) );
  AOI22_X1 U2384 ( .A1(n2442), .A2(\xmem_inst/mem[3][7] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][7] ), .ZN(n2262) );
  AOI22_X1 U2385 ( .A1(n2885), .A2(\xmem_inst/mem[2][7] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][7] ), .ZN(n2261) );
  NAND4_X1 U2386 ( .A1(n2264), .A2(n2263), .A3(n2262), .A4(n2261), .ZN(n2273)
         );
  AOI22_X1 U2387 ( .A1(n2200), .A2(\xmem_inst/mem[8][7] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][7] ), .ZN(n2268) );
  AOI22_X1 U2388 ( .A1(n2202), .A2(\xmem_inst/mem[14][7] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][7] ), .ZN(n2267) );
  AOI22_X1 U2389 ( .A1(n2447), .A2(\xmem_inst/mem[19][7] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][7] ), .ZN(n2266) );
  AOI22_X1 U2390 ( .A1(n2205), .A2(\xmem_inst/mem[6][7] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][7] ), .ZN(n2265) );
  NAND4_X1 U2391 ( .A1(n2268), .A2(n2267), .A3(n2266), .A4(n2265), .ZN(n2272)
         );
  AOI22_X1 U2392 ( .A1(n3207), .A2(\xmem_inst/mem[16][7] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][7] ), .ZN(n2270) );
  AOI22_X1 U2393 ( .A1(n2214), .A2(\xmem_inst/mem[10][7] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][7] ), .ZN(n2269) );
  NAND2_X1 U2394 ( .A1(n2270), .A2(n2269), .ZN(n2271) );
  AOI22_X1 U2395 ( .A1(n2835), .A2(\xmem_inst/mem[15][1] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][1] ), .ZN(n2277) );
  AOI22_X1 U2396 ( .A1(n2575), .A2(\xmem_inst/mem[7][1] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][1] ), .ZN(n2276) );
  AOI22_X1 U2397 ( .A1(n2442), .A2(\xmem_inst/mem[3][1] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][1] ), .ZN(n2275) );
  AOI22_X1 U2398 ( .A1(n2885), .A2(\xmem_inst/mem[2][1] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][1] ), .ZN(n2274) );
  NAND4_X1 U2399 ( .A1(n2277), .A2(n2276), .A3(n2275), .A4(n2274), .ZN(n2286)
         );
  AOI22_X1 U2400 ( .A1(n2200), .A2(\xmem_inst/mem[8][1] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][1] ), .ZN(n2281) );
  AOI22_X1 U2401 ( .A1(n2202), .A2(\xmem_inst/mem[14][1] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][1] ), .ZN(n2280) );
  AOI22_X1 U2402 ( .A1(n2447), .A2(\xmem_inst/mem[19][1] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][1] ), .ZN(n2279) );
  AOI22_X1 U2403 ( .A1(n2205), .A2(\xmem_inst/mem[6][1] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][1] ), .ZN(n2278) );
  NAND4_X1 U2404 ( .A1(n2281), .A2(n2280), .A3(n2279), .A4(n2278), .ZN(n2285)
         );
  AOI22_X1 U2405 ( .A1(n3207), .A2(\xmem_inst/mem[16][1] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][1] ), .ZN(n2283) );
  AOI22_X1 U2406 ( .A1(n2214), .A2(\xmem_inst/mem[10][1] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][1] ), .ZN(n2282) );
  NAND2_X1 U2407 ( .A1(n2283), .A2(n2282), .ZN(n2284) );
  BUF_X2 U2408 ( .A(n2287), .Z(n2379) );
  AND2_X1 U2409 ( .A1(n2291), .A2(n2319), .ZN(n2288) );
  INV_X1 U2410 ( .A(n2294), .ZN(n2383) );
  NAND2_X1 U2411 ( .A1(n2383), .A2(n2375), .ZN(n2295) );
  XNOR2_X1 U2412 ( .A(n2391), .B(n2295), .ZN(n2296) );
  NAND2_X1 U2413 ( .A1(n2379), .A2(n2296), .ZN(n2297) );
  NAND3_X1 U2414 ( .A1(n2297), .A2(n2399), .A3(n1362), .ZN(n894) );
  AND2_X1 U2415 ( .A1(\DP_OP_485J1_122_4413/n1204 ), .A2(xmem_data[0]), .ZN(
        n2298) );
  NAND2_X1 U2416 ( .A1(n2397), .A2(n2298), .ZN(n2299) );
  NAND3_X1 U2417 ( .A1(n2299), .A2(n2399), .A3(n1363), .ZN(n910) );
  OR2_X1 U2418 ( .A1(n2301), .A2(n2300), .ZN(n2303) );
  AND2_X1 U2419 ( .A1(n2303), .A2(n2302), .ZN(n2304) );
  NAND2_X1 U2420 ( .A1(n2397), .A2(n2304), .ZN(n2305) );
  NAND3_X1 U2421 ( .A1(n2305), .A2(n2399), .A3(n1364), .ZN(n909) );
  NAND2_X1 U2422 ( .A1(n2307), .A2(n2306), .ZN(n2309) );
  XNOR2_X1 U2423 ( .A(n2309), .B(n2308), .ZN(n2310) );
  NAND2_X1 U2424 ( .A1(n2379), .A2(n2310), .ZN(n2311) );
  NAND3_X1 U2425 ( .A1(n2311), .A2(n2399), .A3(n1365), .ZN(n908) );
  OAI21_X1 U2426 ( .B1(n2323), .B2(n2175), .A(n2312), .ZN(n2316) );
  NAND2_X1 U2427 ( .A1(n2314), .A2(n2313), .ZN(n2315) );
  XNOR2_X1 U2428 ( .A(n2316), .B(n2315), .ZN(n2317) );
  NAND2_X1 U2429 ( .A1(n2379), .A2(n2317), .ZN(n2318) );
  NAND3_X1 U2430 ( .A1(n2318), .A2(n2399), .A3(n1366), .ZN(n897) );
  INV_X1 U2431 ( .A(n2319), .ZN(n2322) );
  INV_X1 U2432 ( .A(n2320), .ZN(n2321) );
  OAI21_X1 U2433 ( .B1(n2323), .B2(n2322), .A(n2321), .ZN(n2328) );
  INV_X1 U2434 ( .A(n2324), .ZN(n2326) );
  NAND2_X1 U2435 ( .A1(n2326), .A2(n2325), .ZN(n2327) );
  XNOR2_X1 U2436 ( .A(n2328), .B(n2327), .ZN(n2329) );
  NAND2_X1 U2437 ( .A1(n2379), .A2(n2329), .ZN(n2330) );
  NAND2_X2 U2438 ( .A1(n2794), .A2(n2796), .ZN(n2381) );
  NAND3_X1 U2439 ( .A1(n2330), .A2(n2381), .A3(n1367), .ZN(n896) );
  INV_X1 U2440 ( .A(n2331), .ZN(n2333) );
  NAND2_X1 U2441 ( .A1(n2333), .A2(n2332), .ZN(n2335) );
  XOR2_X1 U2442 ( .A(n2335), .B(n2334), .Z(n2336) );
  NAND2_X1 U2443 ( .A1(n2379), .A2(n2336), .ZN(n2337) );
  NAND3_X1 U2444 ( .A1(n2337), .A2(n2381), .A3(n1368), .ZN(n907) );
  INV_X1 U2445 ( .A(n2338), .ZN(n2340) );
  NAND2_X1 U2446 ( .A1(n2340), .A2(n2339), .ZN(n2341) );
  XOR2_X1 U2447 ( .A(n2342), .B(n2341), .Z(n2343) );
  NAND2_X1 U2448 ( .A1(n2379), .A2(n2343), .ZN(n2344) );
  NAND3_X1 U2449 ( .A1(n2344), .A2(n2381), .A3(n1369), .ZN(n905) );
  INV_X1 U2450 ( .A(n2346), .ZN(n2347) );
  AOI21_X1 U2451 ( .B1(n2191), .B2(n2348), .A(n2347), .ZN(n2352) );
  NAND2_X1 U2452 ( .A1(n2350), .A2(n2349), .ZN(n2351) );
  XOR2_X1 U2453 ( .A(n2352), .B(n2351), .Z(n2353) );
  NAND2_X1 U2454 ( .A1(n2379), .A2(n2353), .ZN(n2354) );
  NAND3_X1 U2455 ( .A1(n2354), .A2(n2381), .A3(n1370), .ZN(n899) );
  NAND2_X1 U2456 ( .A1(n2356), .A2(n2355), .ZN(n2357) );
  XOR2_X1 U2457 ( .A(n2358), .B(n2357), .Z(n2359) );
  NAND2_X1 U2458 ( .A1(n2379), .A2(n2359), .ZN(n2360) );
  NAND3_X1 U2459 ( .A1(n2360), .A2(n2381), .A3(n1371), .ZN(n903) );
  NAND2_X1 U2460 ( .A1(n2362), .A2(n2361), .ZN(n2363) );
  XOR2_X1 U2461 ( .A(n2364), .B(n2363), .Z(n2365) );
  NAND2_X1 U2462 ( .A1(n2379), .A2(n2365), .ZN(n2366) );
  NAND3_X1 U2463 ( .A1(n2366), .A2(n2381), .A3(n1372), .ZN(n901) );
  INV_X1 U2464 ( .A(n2368), .ZN(n2370) );
  AND2_X1 U2465 ( .A1(n2370), .A2(n2369), .ZN(n2371) );
  XNOR2_X1 U2466 ( .A(n2372), .B(n2371), .ZN(n2373) );
  NAND2_X1 U2467 ( .A1(n2379), .A2(n2373), .ZN(n2374) );
  NAND3_X1 U2468 ( .A1(n2374), .A2(n2381), .A3(n1373), .ZN(n895) );
  INV_X1 U2469 ( .A(n2375), .ZN(n2386) );
  AOI21_X1 U2470 ( .B1(n2391), .B2(n2383), .A(n2386), .ZN(n2378) );
  INV_X1 U2471 ( .A(n1344), .ZN(n2387) );
  AND2_X1 U2472 ( .A1(n2387), .A2(n2384), .ZN(n2377) );
  XNOR2_X1 U2473 ( .A(n2378), .B(n2377), .ZN(n2380) );
  NAND2_X1 U2474 ( .A1(n2380), .A2(n2379), .ZN(n2382) );
  NAND3_X1 U2475 ( .A1(n2382), .A2(n2381), .A3(n1374), .ZN(n893) );
  AND2_X1 U2476 ( .A1(n2383), .A2(n2387), .ZN(n2390) );
  INV_X1 U2477 ( .A(n2384), .ZN(n2385) );
  AOI21_X1 U2478 ( .B1(n2387), .B2(n2386), .A(n2385), .ZN(n2388) );
  INV_X1 U2479 ( .A(n2388), .ZN(n2389) );
  AOI21_X1 U2480 ( .B1(n2391), .B2(n2390), .A(n2389), .ZN(n2396) );
  INV_X1 U2481 ( .A(n2392), .ZN(n2394) );
  AND2_X1 U2482 ( .A1(n2394), .A2(n2393), .ZN(n2395) );
  XNOR2_X1 U2483 ( .A(n2396), .B(n2395), .ZN(n2398) );
  NAND2_X1 U2484 ( .A1(n2398), .A2(n2397), .ZN(n2400) );
  NAND3_X1 U2485 ( .A1(n2400), .A2(n2399), .A3(n1375), .ZN(n892) );
  AOI22_X1 U2486 ( .A1(\xmem_inst/mem[10][0] ), .A2(n2214), .B1(
        \xmem_inst/mem[12][0] ), .B2(n2216), .ZN(n2402) );
  AOI22_X1 U2487 ( .A1(\xmem_inst/mem[14][0] ), .A2(n2202), .B1(
        \xmem_inst/mem[11][0] ), .B2(n2203), .ZN(n2401) );
  NAND2_X1 U2488 ( .A1(n2402), .A2(n2401), .ZN(n2414) );
  AOI22_X1 U2489 ( .A1(n2835), .A2(\xmem_inst/mem[15][0] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][0] ), .ZN(n2405) );
  AOI22_X1 U2490 ( .A1(n2885), .A2(\xmem_inst/mem[2][0] ), .B1(n2442), .B2(
        \xmem_inst/mem[3][0] ), .ZN(n2404) );
  AOI22_X1 U2491 ( .A1(n2415), .A2(\xmem_inst/mem[0][0] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][0] ), .ZN(n2403) );
  NAND3_X1 U2492 ( .A1(n2405), .A2(n2404), .A3(n2403), .ZN(n2413) );
  AOI22_X1 U2493 ( .A1(\xmem_inst/mem[8][0] ), .A2(n2200), .B1(
        \xmem_inst/mem[5][0] ), .B2(n2201), .ZN(n2407) );
  AOI22_X1 U2494 ( .A1(\xmem_inst/mem[6][0] ), .A2(n2205), .B1(
        \xmem_inst/mem[4][0] ), .B2(n2207), .ZN(n2406) );
  NAND2_X1 U2495 ( .A1(n2407), .A2(n2406), .ZN(n2412) );
  AOI22_X1 U2496 ( .A1(\xmem_inst/mem[13][0] ), .A2(n2212), .B1(n2204), .B2(
        \xmem_inst/mem[9][0] ), .ZN(n2410) );
  AOI22_X1 U2497 ( .A1(n2575), .A2(\xmem_inst/mem[7][0] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][0] ), .ZN(n2409) );
  AOI22_X1 U2498 ( .A1(n3207), .A2(\xmem_inst/mem[16][0] ), .B1(
        \xmem_inst/mem[19][0] ), .B2(n2447), .ZN(n2408) );
  NAND3_X1 U2499 ( .A1(n2410), .A2(n2409), .A3(n2408), .ZN(n2411) );
  OR4_X1 U2500 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .ZN(
        \xmem_inst/N109 ) );
  AOI22_X1 U2501 ( .A1(n2835), .A2(\xmem_inst/mem[15][9] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][9] ), .ZN(n2419) );
  AOI22_X1 U2502 ( .A1(n2575), .A2(\xmem_inst/mem[7][9] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][9] ), .ZN(n2418) );
  AOI22_X1 U2503 ( .A1(n2442), .A2(\xmem_inst/mem[3][9] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][9] ), .ZN(n2417) );
  AOI22_X1 U2504 ( .A1(n2885), .A2(\xmem_inst/mem[2][9] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][9] ), .ZN(n2416) );
  NAND4_X1 U2505 ( .A1(n2419), .A2(n2418), .A3(n2417), .A4(n2416), .ZN(n2428)
         );
  AOI22_X1 U2506 ( .A1(n2200), .A2(\xmem_inst/mem[8][9] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][9] ), .ZN(n2423) );
  AOI22_X1 U2507 ( .A1(n2202), .A2(\xmem_inst/mem[14][9] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][9] ), .ZN(n2422) );
  AOI22_X1 U2508 ( .A1(n2447), .A2(\xmem_inst/mem[19][9] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][9] ), .ZN(n2421) );
  AOI22_X1 U2509 ( .A1(n2205), .A2(\xmem_inst/mem[6][9] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][9] ), .ZN(n2420) );
  NAND4_X1 U2510 ( .A1(n2423), .A2(n2422), .A3(n2421), .A4(n2420), .ZN(n2427)
         );
  AOI22_X1 U2511 ( .A1(n3207), .A2(\xmem_inst/mem[16][9] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][9] ), .ZN(n2425) );
  AOI22_X1 U2512 ( .A1(n2214), .A2(\xmem_inst/mem[10][9] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][9] ), .ZN(n2424) );
  NAND2_X1 U2513 ( .A1(n2425), .A2(n2424), .ZN(n2426) );
  OR3_X1 U2514 ( .A1(n2428), .A2(n2427), .A3(n2426), .ZN(\xmem_inst/N100 ) );
  AOI22_X1 U2515 ( .A1(n2835), .A2(\xmem_inst/mem[15][10] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][10] ), .ZN(n2432) );
  AOI22_X1 U2516 ( .A1(n2575), .A2(\xmem_inst/mem[7][10] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][10] ), .ZN(n2431) );
  AOI22_X1 U2517 ( .A1(n2442), .A2(\xmem_inst/mem[3][10] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][10] ), .ZN(n2430) );
  AOI22_X1 U2518 ( .A1(n2885), .A2(\xmem_inst/mem[2][10] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][10] ), .ZN(n2429) );
  NAND4_X1 U2519 ( .A1(n2432), .A2(n2431), .A3(n2430), .A4(n2429), .ZN(n2441)
         );
  AOI22_X1 U2520 ( .A1(n2200), .A2(\xmem_inst/mem[8][10] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][10] ), .ZN(n2436) );
  AOI22_X1 U2521 ( .A1(n2202), .A2(\xmem_inst/mem[14][10] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][10] ), .ZN(n2435) );
  AOI22_X1 U2522 ( .A1(n2447), .A2(\xmem_inst/mem[19][10] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][10] ), .ZN(n2434) );
  AOI22_X1 U2523 ( .A1(n2205), .A2(\xmem_inst/mem[6][10] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][10] ), .ZN(n2433) );
  NAND4_X1 U2524 ( .A1(n2436), .A2(n2435), .A3(n2434), .A4(n2433), .ZN(n2440)
         );
  AOI22_X1 U2525 ( .A1(n3207), .A2(\xmem_inst/mem[16][10] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][10] ), .ZN(n2438) );
  AOI22_X1 U2526 ( .A1(n2214), .A2(\xmem_inst/mem[10][10] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][10] ), .ZN(n2437) );
  NAND2_X1 U2527 ( .A1(n2438), .A2(n2437), .ZN(n2439) );
  OR3_X1 U2528 ( .A1(n2441), .A2(n2440), .A3(n2439), .ZN(\xmem_inst/N99 ) );
  AOI22_X1 U2529 ( .A1(n2835), .A2(\xmem_inst/mem[15][2] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][2] ), .ZN(n2446) );
  AOI22_X1 U2530 ( .A1(n2575), .A2(\xmem_inst/mem[7][2] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][2] ), .ZN(n2445) );
  AOI22_X1 U2531 ( .A1(n2442), .A2(\xmem_inst/mem[3][2] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][2] ), .ZN(n2444) );
  AOI22_X1 U2532 ( .A1(n2885), .A2(\xmem_inst/mem[2][2] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][2] ), .ZN(n2443) );
  NAND4_X1 U2533 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n2456)
         );
  AOI22_X1 U2534 ( .A1(n2200), .A2(\xmem_inst/mem[8][2] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][2] ), .ZN(n2451) );
  AOI22_X1 U2535 ( .A1(n2202), .A2(\xmem_inst/mem[14][2] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][2] ), .ZN(n2450) );
  AOI22_X1 U2536 ( .A1(n2447), .A2(\xmem_inst/mem[19][2] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][2] ), .ZN(n2449) );
  AOI22_X1 U2537 ( .A1(n2205), .A2(\xmem_inst/mem[6][2] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][2] ), .ZN(n2448) );
  NAND4_X1 U2538 ( .A1(n2451), .A2(n2450), .A3(n2449), .A4(n2448), .ZN(n2455)
         );
  AOI22_X1 U2539 ( .A1(n3207), .A2(\xmem_inst/mem[16][2] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][2] ), .ZN(n2453) );
  AOI22_X1 U2540 ( .A1(n2214), .A2(\xmem_inst/mem[10][2] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][2] ), .ZN(n2452) );
  NAND2_X1 U2541 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  OR3_X1 U2542 ( .A1(n2456), .A2(n2455), .A3(n2454), .ZN(\xmem_inst/N107 ) );
  AOI22_X1 U2543 ( .A1(n2835), .A2(\xmem_inst/mem[15][6] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][6] ), .ZN(n2461) );
  AOI22_X1 U2544 ( .A1(n2575), .A2(\xmem_inst/mem[7][6] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][6] ), .ZN(n2460) );
  AOI22_X1 U2545 ( .A1(n2442), .A2(\xmem_inst/mem[3][6] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][6] ), .ZN(n2459) );
  AOI22_X1 U2546 ( .A1(n2885), .A2(\xmem_inst/mem[2][6] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][6] ), .ZN(n2458) );
  NAND4_X1 U2547 ( .A1(n2461), .A2(n2460), .A3(n2459), .A4(n2458), .ZN(n2470)
         );
  AOI22_X1 U2548 ( .A1(n2200), .A2(\xmem_inst/mem[8][6] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][6] ), .ZN(n2465) );
  AOI22_X1 U2549 ( .A1(n2202), .A2(\xmem_inst/mem[14][6] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][6] ), .ZN(n2464) );
  AOI22_X1 U2550 ( .A1(n2447), .A2(\xmem_inst/mem[19][6] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][6] ), .ZN(n2463) );
  AOI22_X1 U2551 ( .A1(n2205), .A2(\xmem_inst/mem[6][6] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][6] ), .ZN(n2462) );
  NAND4_X1 U2552 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n2469)
         );
  AOI22_X1 U2553 ( .A1(n3207), .A2(\xmem_inst/mem[16][6] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][6] ), .ZN(n2467) );
  AOI22_X1 U2554 ( .A1(n2214), .A2(\xmem_inst/mem[10][6] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][6] ), .ZN(n2466) );
  NAND2_X1 U2555 ( .A1(n2467), .A2(n2466), .ZN(n2468) );
  OR3_X1 U2556 ( .A1(n2470), .A2(n2469), .A3(n2468), .ZN(\xmem_inst/N103 ) );
  AOI22_X1 U2557 ( .A1(n2835), .A2(\xmem_inst/mem[15][15] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][15] ), .ZN(n2474) );
  AOI22_X1 U2558 ( .A1(n2575), .A2(\xmem_inst/mem[7][15] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][15] ), .ZN(n2473) );
  AOI22_X1 U2559 ( .A1(n2442), .A2(\xmem_inst/mem[3][15] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][15] ), .ZN(n2472) );
  AOI22_X1 U2560 ( .A1(n2885), .A2(\xmem_inst/mem[2][15] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][15] ), .ZN(n2471) );
  NAND4_X1 U2561 ( .A1(n2474), .A2(n2473), .A3(n2472), .A4(n2471), .ZN(n2483)
         );
  AOI22_X1 U2562 ( .A1(n2200), .A2(\xmem_inst/mem[8][15] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][15] ), .ZN(n2478) );
  AOI22_X1 U2563 ( .A1(n2202), .A2(\xmem_inst/mem[14][15] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][15] ), .ZN(n2477) );
  AOI22_X1 U2564 ( .A1(n2447), .A2(\xmem_inst/mem[19][15] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][15] ), .ZN(n2476) );
  AOI22_X1 U2565 ( .A1(n2205), .A2(\xmem_inst/mem[6][15] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][15] ), .ZN(n2475) );
  NAND4_X1 U2566 ( .A1(n2478), .A2(n2477), .A3(n2476), .A4(n2475), .ZN(n2482)
         );
  AOI22_X1 U2567 ( .A1(n3207), .A2(\xmem_inst/mem[16][15] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][15] ), .ZN(n2480) );
  AOI22_X1 U2568 ( .A1(n2214), .A2(\xmem_inst/mem[10][15] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][15] ), .ZN(n2479) );
  NAND2_X1 U2569 ( .A1(n2480), .A2(n2479), .ZN(n2481) );
  OR3_X1 U2570 ( .A1(n2483), .A2(n2482), .A3(n2481), .ZN(\xmem_inst/N94 ) );
  AOI22_X1 U2571 ( .A1(n2835), .A2(\xmem_inst/mem[15][11] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][11] ), .ZN(n2487) );
  AOI22_X1 U2572 ( .A1(n2575), .A2(\xmem_inst/mem[7][11] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][11] ), .ZN(n2486) );
  AOI22_X1 U2573 ( .A1(n2442), .A2(\xmem_inst/mem[3][11] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][11] ), .ZN(n2485) );
  AOI22_X1 U2574 ( .A1(n2885), .A2(\xmem_inst/mem[2][11] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][11] ), .ZN(n2484) );
  NAND4_X1 U2575 ( .A1(n2487), .A2(n2486), .A3(n2485), .A4(n2484), .ZN(n2496)
         );
  AOI22_X1 U2576 ( .A1(n2200), .A2(\xmem_inst/mem[8][11] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][11] ), .ZN(n2491) );
  AOI22_X1 U2577 ( .A1(n2202), .A2(\xmem_inst/mem[14][11] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][11] ), .ZN(n2490) );
  AOI22_X1 U2578 ( .A1(n2447), .A2(\xmem_inst/mem[19][11] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][11] ), .ZN(n2489) );
  AOI22_X1 U2579 ( .A1(n2205), .A2(\xmem_inst/mem[6][11] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][11] ), .ZN(n2488) );
  NAND4_X1 U2580 ( .A1(n2491), .A2(n2490), .A3(n2489), .A4(n2488), .ZN(n2495)
         );
  AOI22_X1 U2581 ( .A1(n3207), .A2(\xmem_inst/mem[16][11] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][11] ), .ZN(n2493) );
  AOI22_X1 U2582 ( .A1(n2214), .A2(\xmem_inst/mem[10][11] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][11] ), .ZN(n2492) );
  NAND2_X1 U2583 ( .A1(n2493), .A2(n2492), .ZN(n2494) );
  OR3_X1 U2584 ( .A1(n2496), .A2(n2495), .A3(n2494), .ZN(\xmem_inst/N98 ) );
  AOI22_X1 U2585 ( .A1(n2835), .A2(\xmem_inst/mem[15][3] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][3] ), .ZN(n2500) );
  AOI22_X1 U2586 ( .A1(n2575), .A2(\xmem_inst/mem[7][3] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][3] ), .ZN(n2499) );
  AOI22_X1 U2587 ( .A1(n2442), .A2(\xmem_inst/mem[3][3] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][3] ), .ZN(n2498) );
  AOI22_X1 U2588 ( .A1(n2885), .A2(\xmem_inst/mem[2][3] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][3] ), .ZN(n2497) );
  NAND4_X1 U2589 ( .A1(n2500), .A2(n2499), .A3(n2498), .A4(n2497), .ZN(n2509)
         );
  AOI22_X1 U2590 ( .A1(n2200), .A2(\xmem_inst/mem[8][3] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][3] ), .ZN(n2504) );
  AOI22_X1 U2591 ( .A1(n2202), .A2(\xmem_inst/mem[14][3] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][3] ), .ZN(n2503) );
  AOI22_X1 U2592 ( .A1(n2447), .A2(\xmem_inst/mem[19][3] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][3] ), .ZN(n2502) );
  AOI22_X1 U2593 ( .A1(n2205), .A2(\xmem_inst/mem[6][3] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][3] ), .ZN(n2501) );
  NAND4_X1 U2594 ( .A1(n2504), .A2(n2503), .A3(n2502), .A4(n2501), .ZN(n2508)
         );
  AOI22_X1 U2595 ( .A1(n3207), .A2(\xmem_inst/mem[16][3] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][3] ), .ZN(n2506) );
  AOI22_X1 U2596 ( .A1(n2214), .A2(\xmem_inst/mem[10][3] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][3] ), .ZN(n2505) );
  NAND2_X1 U2597 ( .A1(n2506), .A2(n2505), .ZN(n2507) );
  OR3_X1 U2598 ( .A1(n2509), .A2(n2508), .A3(n2507), .ZN(\xmem_inst/N106 ) );
  AOI22_X1 U2599 ( .A1(n2835), .A2(\xmem_inst/mem[15][4] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][4] ), .ZN(n2513) );
  AOI22_X1 U2600 ( .A1(n2575), .A2(\xmem_inst/mem[7][4] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][4] ), .ZN(n2512) );
  AOI22_X1 U2601 ( .A1(n2442), .A2(\xmem_inst/mem[3][4] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][4] ), .ZN(n2511) );
  AOI22_X1 U2602 ( .A1(n2885), .A2(\xmem_inst/mem[2][4] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][4] ), .ZN(n2510) );
  NAND4_X1 U2603 ( .A1(n2513), .A2(n2512), .A3(n2511), .A4(n2510), .ZN(n2522)
         );
  AOI22_X1 U2604 ( .A1(n2200), .A2(\xmem_inst/mem[8][4] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][4] ), .ZN(n2517) );
  AOI22_X1 U2605 ( .A1(n2202), .A2(\xmem_inst/mem[14][4] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][4] ), .ZN(n2516) );
  AOI22_X1 U2606 ( .A1(n2447), .A2(\xmem_inst/mem[19][4] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][4] ), .ZN(n2515) );
  AOI22_X1 U2607 ( .A1(n2205), .A2(\xmem_inst/mem[6][4] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][4] ), .ZN(n2514) );
  NAND4_X1 U2608 ( .A1(n2517), .A2(n2516), .A3(n2515), .A4(n2514), .ZN(n2521)
         );
  AOI22_X1 U2609 ( .A1(n3207), .A2(\xmem_inst/mem[16][4] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][4] ), .ZN(n2519) );
  AOI22_X1 U2610 ( .A1(n2214), .A2(\xmem_inst/mem[10][4] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][4] ), .ZN(n2518) );
  NAND2_X1 U2611 ( .A1(n2519), .A2(n2518), .ZN(n2520) );
  OR3_X1 U2612 ( .A1(n2522), .A2(n2521), .A3(n2520), .ZN(\xmem_inst/N105 ) );
  AOI22_X1 U2613 ( .A1(n2835), .A2(\xmem_inst/mem[15][8] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][8] ), .ZN(n2526) );
  AOI22_X1 U2614 ( .A1(n2575), .A2(\xmem_inst/mem[7][8] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][8] ), .ZN(n2525) );
  AOI22_X1 U2615 ( .A1(n2442), .A2(\xmem_inst/mem[3][8] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][8] ), .ZN(n2524) );
  AOI22_X1 U2616 ( .A1(n2885), .A2(\xmem_inst/mem[2][8] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][8] ), .ZN(n2523) );
  NAND4_X1 U2617 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n2535)
         );
  AOI22_X1 U2618 ( .A1(n2200), .A2(\xmem_inst/mem[8][8] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][8] ), .ZN(n2530) );
  AOI22_X1 U2619 ( .A1(n2202), .A2(\xmem_inst/mem[14][8] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][8] ), .ZN(n2529) );
  AOI22_X1 U2620 ( .A1(n2447), .A2(\xmem_inst/mem[19][8] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][8] ), .ZN(n2528) );
  AOI22_X1 U2621 ( .A1(n2205), .A2(\xmem_inst/mem[6][8] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][8] ), .ZN(n2527) );
  NAND4_X1 U2622 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n2534)
         );
  AOI22_X1 U2623 ( .A1(n3207), .A2(\xmem_inst/mem[16][8] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][8] ), .ZN(n2532) );
  AOI22_X1 U2624 ( .A1(n2214), .A2(\xmem_inst/mem[10][8] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][8] ), .ZN(n2531) );
  NAND2_X1 U2625 ( .A1(n2532), .A2(n2531), .ZN(n2533) );
  OR3_X1 U2626 ( .A1(n2535), .A2(n2534), .A3(n2533), .ZN(\xmem_inst/N101 ) );
  AOI22_X1 U2627 ( .A1(n2835), .A2(\xmem_inst/mem[15][18] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][18] ), .ZN(n2539) );
  AOI22_X1 U2628 ( .A1(n2575), .A2(\xmem_inst/mem[7][18] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][18] ), .ZN(n2538) );
  AOI22_X1 U2629 ( .A1(n2442), .A2(\xmem_inst/mem[3][18] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][18] ), .ZN(n2537) );
  AOI22_X1 U2630 ( .A1(n2885), .A2(\xmem_inst/mem[2][18] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][18] ), .ZN(n2536) );
  NAND4_X1 U2631 ( .A1(n2539), .A2(n2538), .A3(n2537), .A4(n2536), .ZN(n2548)
         );
  AOI22_X1 U2632 ( .A1(n2200), .A2(\xmem_inst/mem[8][18] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][18] ), .ZN(n2543) );
  AOI22_X1 U2633 ( .A1(n2202), .A2(\xmem_inst/mem[14][18] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][18] ), .ZN(n2542) );
  AOI22_X1 U2634 ( .A1(n2447), .A2(\xmem_inst/mem[19][18] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][18] ), .ZN(n2541) );
  AOI22_X1 U2635 ( .A1(n2205), .A2(\xmem_inst/mem[6][18] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][18] ), .ZN(n2540) );
  NAND4_X1 U2636 ( .A1(n2543), .A2(n2542), .A3(n2541), .A4(n2540), .ZN(n2547)
         );
  AOI22_X1 U2637 ( .A1(n3207), .A2(\xmem_inst/mem[16][18] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][18] ), .ZN(n2545) );
  AOI22_X1 U2638 ( .A1(n2214), .A2(\xmem_inst/mem[10][18] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][18] ), .ZN(n2544) );
  NAND2_X1 U2639 ( .A1(n2545), .A2(n2544), .ZN(n2546) );
  OR3_X1 U2640 ( .A1(n2548), .A2(n2547), .A3(n2546), .ZN(\xmem_inst/N91 ) );
  AOI22_X1 U2641 ( .A1(n2835), .A2(\xmem_inst/mem[15][12] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][12] ), .ZN(n2552) );
  AOI22_X1 U2642 ( .A1(n2575), .A2(\xmem_inst/mem[7][12] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][12] ), .ZN(n2551) );
  AOI22_X1 U2643 ( .A1(n2442), .A2(\xmem_inst/mem[3][12] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][12] ), .ZN(n2550) );
  AOI22_X1 U2644 ( .A1(n2885), .A2(\xmem_inst/mem[2][12] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][12] ), .ZN(n2549) );
  NAND4_X1 U2645 ( .A1(n2552), .A2(n2551), .A3(n2550), .A4(n2549), .ZN(n2561)
         );
  AOI22_X1 U2646 ( .A1(n2200), .A2(\xmem_inst/mem[8][12] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][12] ), .ZN(n2556) );
  AOI22_X1 U2647 ( .A1(n2202), .A2(\xmem_inst/mem[14][12] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][12] ), .ZN(n2555) );
  AOI22_X1 U2648 ( .A1(n2447), .A2(\xmem_inst/mem[19][12] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][12] ), .ZN(n2554) );
  AOI22_X1 U2649 ( .A1(n2205), .A2(\xmem_inst/mem[6][12] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][12] ), .ZN(n2553) );
  NAND4_X1 U2650 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n2560)
         );
  AOI22_X1 U2651 ( .A1(n3207), .A2(\xmem_inst/mem[16][12] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][12] ), .ZN(n2558) );
  AOI22_X1 U2652 ( .A1(n2214), .A2(\xmem_inst/mem[10][12] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][12] ), .ZN(n2557) );
  NAND2_X1 U2653 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  OR3_X1 U2654 ( .A1(n2561), .A2(n2560), .A3(n2559), .ZN(\xmem_inst/N97 ) );
  AOI22_X1 U2655 ( .A1(n2835), .A2(\xmem_inst/mem[15][16] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][16] ), .ZN(n2565) );
  AOI22_X1 U2656 ( .A1(n2575), .A2(\xmem_inst/mem[7][16] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][16] ), .ZN(n2564) );
  AOI22_X1 U2657 ( .A1(n2442), .A2(\xmem_inst/mem[3][16] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][16] ), .ZN(n2563) );
  AOI22_X1 U2658 ( .A1(n2885), .A2(\xmem_inst/mem[2][16] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][16] ), .ZN(n2562) );
  NAND4_X1 U2659 ( .A1(n2565), .A2(n2564), .A3(n2563), .A4(n2562), .ZN(n2574)
         );
  AOI22_X1 U2660 ( .A1(n2200), .A2(\xmem_inst/mem[8][16] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][16] ), .ZN(n2569) );
  AOI22_X1 U2661 ( .A1(n2202), .A2(\xmem_inst/mem[14][16] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][16] ), .ZN(n2568) );
  AOI22_X1 U2662 ( .A1(n2447), .A2(\xmem_inst/mem[19][16] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][16] ), .ZN(n2567) );
  AOI22_X1 U2663 ( .A1(n2205), .A2(\xmem_inst/mem[6][16] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][16] ), .ZN(n2566) );
  NAND4_X1 U2664 ( .A1(n2569), .A2(n2568), .A3(n2567), .A4(n2566), .ZN(n2573)
         );
  AOI22_X1 U2665 ( .A1(n3207), .A2(\xmem_inst/mem[16][16] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][16] ), .ZN(n2571) );
  AOI22_X1 U2666 ( .A1(n2214), .A2(\xmem_inst/mem[10][16] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][16] ), .ZN(n2570) );
  NAND2_X1 U2667 ( .A1(n2571), .A2(n2570), .ZN(n2572) );
  OR3_X1 U2668 ( .A1(n2574), .A2(n2573), .A3(n2572), .ZN(\xmem_inst/N93 ) );
  AOI22_X1 U2669 ( .A1(n2835), .A2(\xmem_inst/mem[15][14] ), .B1(n3230), .B2(
        \xmem_inst/mem[17][14] ), .ZN(n2579) );
  AOI22_X1 U2670 ( .A1(n2575), .A2(\xmem_inst/mem[7][14] ), .B1(n3253), .B2(
        \xmem_inst/mem[18][14] ), .ZN(n2578) );
  AOI22_X1 U2671 ( .A1(n2442), .A2(\xmem_inst/mem[3][14] ), .B1(n2457), .B2(
        \xmem_inst/mem[1][14] ), .ZN(n2577) );
  AOI22_X1 U2672 ( .A1(n2885), .A2(\xmem_inst/mem[2][14] ), .B1(n2415), .B2(
        \xmem_inst/mem[0][14] ), .ZN(n2576) );
  NAND4_X1 U2673 ( .A1(n2579), .A2(n2578), .A3(n2577), .A4(n2576), .ZN(n2588)
         );
  AOI22_X1 U2674 ( .A1(n2200), .A2(\xmem_inst/mem[8][14] ), .B1(n2201), .B2(
        \xmem_inst/mem[5][14] ), .ZN(n2583) );
  AOI22_X1 U2675 ( .A1(n2202), .A2(\xmem_inst/mem[14][14] ), .B1(n2203), .B2(
        \xmem_inst/mem[11][14] ), .ZN(n2582) );
  AOI22_X1 U2676 ( .A1(n2447), .A2(\xmem_inst/mem[19][14] ), .B1(n2204), .B2(
        \xmem_inst/mem[9][14] ), .ZN(n2581) );
  AOI22_X1 U2677 ( .A1(n2205), .A2(\xmem_inst/mem[6][14] ), .B1(n2207), .B2(
        \xmem_inst/mem[4][14] ), .ZN(n2580) );
  NAND4_X1 U2678 ( .A1(n2583), .A2(n2582), .A3(n2581), .A4(n2580), .ZN(n2587)
         );
  AOI22_X1 U2679 ( .A1(n3207), .A2(\xmem_inst/mem[16][14] ), .B1(n2212), .B2(
        \xmem_inst/mem[13][14] ), .ZN(n2585) );
  AOI22_X1 U2680 ( .A1(n2214), .A2(\xmem_inst/mem[10][14] ), .B1(n2216), .B2(
        \xmem_inst/mem[12][14] ), .ZN(n2584) );
  NAND2_X1 U2681 ( .A1(n2585), .A2(n2584), .ZN(n2586) );
  OR3_X1 U2682 ( .A1(n2588), .A2(n2587), .A3(n2586), .ZN(\xmem_inst/N95 ) );
  NAND2_X1 U2683 ( .A1(fmem_addr[2]), .A2(fmem_addr[3]), .ZN(n2639) );
  INV_X1 U2684 ( .A(n2639), .ZN(n2605) );
  NAND2_X1 U2685 ( .A1(n3347), .A2(n3331), .ZN(n2604) );
  NAND2_X1 U2686 ( .A1(n2605), .A2(n2604), .ZN(n2612) );
  NAND2_X1 U2687 ( .A1(n3332), .A2(fmem_addr[3]), .ZN(n3302) );
  INV_X1 U2688 ( .A(n3302), .ZN(n2602) );
  NAND2_X1 U2689 ( .A1(fmem_addr[0]), .A2(fmem_addr[1]), .ZN(n2640) );
  AOI221_X1 U2690 ( .B1(fmem_addr[1]), .B2(fmem_addr[2]), .C1(n3347), .C2(
        n3332), .A(fmem_addr[3]), .ZN(n2601) );
  AOI21_X1 U2691 ( .B1(n2602), .B2(n2640), .A(n2601), .ZN(n2589) );
  OAI21_X1 U2692 ( .B1(n2612), .B2(n3346), .A(n2589), .ZN(n922) );
  NOR2_X1 U2693 ( .A1(fmem_addr[1]), .A2(fmem_addr[3]), .ZN(n2590) );
  NAND2_X1 U2694 ( .A1(n2590), .A2(n3332), .ZN(n2606) );
  OAI211_X1 U2695 ( .C1(n3347), .C2(n3339), .A(fmem_addr[0]), .B(n3332), .ZN(
        n2591) );
  OAI211_X1 U2696 ( .C1(n2612), .C2(n3390), .A(n2606), .B(n2591), .ZN(n918) );
  NAND2_X1 U2697 ( .A1(n3302), .A2(fmem_addr[1]), .ZN(n2592) );
  OAI211_X1 U2698 ( .C1(fmem_addr[1]), .C2(n3339), .A(n2592), .B(n3331), .ZN(
        n2594) );
  XNOR2_X1 U2699 ( .A(fmem_addr[0]), .B(fmem_addr[3]), .ZN(n2593) );
  NAND2_X1 U2700 ( .A1(n2593), .A2(n3332), .ZN(n2613) );
  OAI211_X1 U2701 ( .C1(n2612), .C2(n3389), .A(n2594), .B(n2613), .ZN(n914) );
  NOR3_X1 U2702 ( .A1(fmem_addr[1]), .A2(n3332), .A3(n3331), .ZN(n2596) );
  NOR2_X1 U2703 ( .A1(n3339), .A2(fmem_addr[1]), .ZN(n2610) );
  INV_X1 U2704 ( .A(n2610), .ZN(n2595) );
  OAI22_X1 U2705 ( .A1(n2602), .A2(n2596), .B1(n3331), .B2(n2595), .ZN(n2600)
         );
  OAI211_X1 U2706 ( .C1(n2612), .C2(n1346), .A(n2600), .B(n2606), .ZN(n920) );
  NOR2_X1 U2707 ( .A1(n2639), .A2(n2604), .ZN(n2802) );
  INV_X1 U2708 ( .A(n2802), .ZN(n2597) );
  OAI211_X1 U2709 ( .C1(n2639), .C2(n1347), .A(n2600), .B(n2597), .ZN(n916) );
  NOR2_X1 U2710 ( .A1(fmem_addr[3]), .A2(n3332), .ZN(n2598) );
  NAND2_X1 U2711 ( .A1(n3331), .A2(n2598), .ZN(n2599) );
  OAI211_X1 U2712 ( .C1(n1349), .C2(n2612), .A(n2600), .B(n2599), .ZN(n919) );
  INV_X1 U2713 ( .A(n2640), .ZN(n2603) );
  AOI211_X1 U2714 ( .C1(n2602), .C2(n2603), .A(n2601), .B(n2802), .ZN(n2617)
         );
  NAND3_X1 U2715 ( .A1(n2603), .A2(fmem_addr[2]), .A3(n3339), .ZN(n3306) );
  OAI211_X1 U2716 ( .C1(n2612), .C2(n1348), .A(n2617), .B(n3306), .ZN(n913) );
  NOR2_X1 U2717 ( .A1(n3366), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[18]) );
  NOR2_X1 U2718 ( .A1(n3354), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[6]) );
  NOR2_X1 U2719 ( .A1(n3362), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[15]) );
  NOR2_X1 U2720 ( .A1(n3358), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[10]) );
  NOR2_X1 U2721 ( .A1(n3364), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[11]) );
  NOR2_X1 U2722 ( .A1(n3361), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[14]) );
  NOR2_X1 U2723 ( .A1(n3357), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[9]) );
  NOR2_X1 U2724 ( .A1(n3352), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[4]) );
  NOR2_X1 U2725 ( .A1(n3353), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[5]) );
  NOR2_X1 U2726 ( .A1(n3356), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[8]) );
  NOR2_X1 U2727 ( .A1(n3355), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[7]) );
  NOR2_X1 U2728 ( .A1(n3350), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[2]) );
  NOR2_X1 U2729 ( .A1(n3349), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[1]) );
  NOR2_X1 U2730 ( .A1(n3359), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[12]) );
  INV_X1 U2731 ( .A(n2612), .ZN(n2615) );
  OAI21_X1 U2732 ( .B1(n2605), .B2(n3331), .A(n2604), .ZN(n2607) );
  AOI22_X1 U2733 ( .A1(n2615), .A2(fmem_data[5]), .B1(n2607), .B2(n2606), .ZN(
        n2608) );
  INV_X1 U2734 ( .A(n2608), .ZN(n917) );
  INV_X1 U2735 ( .A(n3306), .ZN(n2609) );
  AOI21_X1 U2736 ( .B1(n2610), .B2(n3331), .A(n2609), .ZN(n2611) );
  OAI211_X1 U2737 ( .C1(n1350), .C2(n2612), .A(n2611), .B(n2613), .ZN(n915) );
  NAND2_X1 U2738 ( .A1(n2615), .A2(fmem_data[1]), .ZN(n2614) );
  OAI211_X1 U2739 ( .C1(fmem_addr[2]), .C2(fmem_addr[1]), .A(n2614), .B(n2613), 
        .ZN(n921) );
  NAND2_X1 U2740 ( .A1(n2615), .A2(fmem_data[19]), .ZN(n2616) );
  OAI211_X1 U2741 ( .C1(fmem_addr[1]), .C2(n3302), .A(n2617), .B(n2616), .ZN(
        n912) );
  NOR2_X1 U2742 ( .A1(n3360), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[13]) );
  NOR2_X1 U2743 ( .A1(n3351), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[3]) );
  NOR2_X1 U2744 ( .A1(n3363), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[16]) );
  NOR2_X1 U2745 ( .A1(n3348), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[0]) );
  NOR2_X1 U2746 ( .A1(n3365), .A2(\mac_unit_inst/adder_reg [19]), .ZN(
        m_data_out_y[17]) );
  NOR2_X1 U2747 ( .A1(n2818), .A2(n3307), .ZN(\ctrl_conv_output_inst/N74 ) );
  NAND2_X1 U2748 ( .A1(m_valid_y), .A2(
        \ctrl_conv_output_inst/conv_start_accum ), .ZN(n2618) );
  NOR2_X1 U2749 ( .A1(\mac_unit_inst/adder_reg [2]), .A2(
        \mac_unit_inst/x_mult_f_reg [2]), .ZN(n2667) );
  NOR2_X1 U2750 ( .A1(\mac_unit_inst/adder_reg [3]), .A2(
        \mac_unit_inst/x_mult_f_reg [3]), .ZN(n2669) );
  NOR2_X1 U2751 ( .A1(n2667), .A2(n2669), .ZN(n2620) );
  NOR2_X1 U2752 ( .A1(\mac_unit_inst/adder_reg [1]), .A2(
        \mac_unit_inst/x_mult_f_reg [1]), .ZN(n2654) );
  NAND2_X1 U2753 ( .A1(\mac_unit_inst/adder_reg [0]), .A2(
        \mac_unit_inst/x_mult_f_reg [0]), .ZN(n2657) );
  NAND2_X1 U2754 ( .A1(\mac_unit_inst/adder_reg [1]), .A2(
        \mac_unit_inst/x_mult_f_reg [1]), .ZN(n2655) );
  OAI21_X1 U2755 ( .B1(n2654), .B2(n2657), .A(n2655), .ZN(n2661) );
  NAND2_X1 U2756 ( .A1(\mac_unit_inst/adder_reg [2]), .A2(
        \mac_unit_inst/x_mult_f_reg [2]), .ZN(n2666) );
  NAND2_X1 U2757 ( .A1(\mac_unit_inst/adder_reg [3]), .A2(
        \mac_unit_inst/x_mult_f_reg [3]), .ZN(n2670) );
  OAI21_X1 U2758 ( .B1(n2669), .B2(n2666), .A(n2670), .ZN(n2619) );
  AOI21_X1 U2759 ( .B1(n2620), .B2(n2661), .A(n2619), .ZN(n2676) );
  NOR2_X1 U2760 ( .A1(\mac_unit_inst/adder_reg [4]), .A2(
        \mac_unit_inst/x_mult_f_reg [4]), .ZN(n2677) );
  NOR2_X1 U2761 ( .A1(\mac_unit_inst/adder_reg [5]), .A2(
        \mac_unit_inst/x_mult_f_reg [5]), .ZN(n2684) );
  NOR2_X1 U2762 ( .A1(n2677), .A2(n2684), .ZN(n2692) );
  NOR2_X1 U2763 ( .A1(\mac_unit_inst/adder_reg [6]), .A2(
        \mac_unit_inst/x_mult_f_reg [6]), .ZN(n2699) );
  NOR2_X1 U2764 ( .A1(\mac_unit_inst/adder_reg [7]), .A2(
        \mac_unit_inst/x_mult_f_reg [7]), .ZN(n2701) );
  NOR2_X1 U2765 ( .A1(n2699), .A2(n2701), .ZN(n2622) );
  NAND2_X1 U2766 ( .A1(n2692), .A2(n2622), .ZN(n2624) );
  NAND2_X1 U2767 ( .A1(\mac_unit_inst/adder_reg [4]), .A2(
        \mac_unit_inst/x_mult_f_reg [4]), .ZN(n2681) );
  NAND2_X1 U2768 ( .A1(\mac_unit_inst/adder_reg [5]), .A2(
        \mac_unit_inst/x_mult_f_reg [5]), .ZN(n2685) );
  OAI21_X1 U2769 ( .B1(n2684), .B2(n2681), .A(n2685), .ZN(n2691) );
  NAND2_X1 U2770 ( .A1(\mac_unit_inst/adder_reg [6]), .A2(
        \mac_unit_inst/x_mult_f_reg [6]), .ZN(n2698) );
  NAND2_X1 U2771 ( .A1(\mac_unit_inst/adder_reg [7]), .A2(
        \mac_unit_inst/x_mult_f_reg [7]), .ZN(n2702) );
  OAI21_X1 U2772 ( .B1(n2701), .B2(n2698), .A(n2702), .ZN(n2621) );
  AOI21_X1 U2773 ( .B1(n2622), .B2(n2691), .A(n2621), .ZN(n2623) );
  OAI21_X1 U2774 ( .B1(n2676), .B2(n2624), .A(n2623), .ZN(n2708) );
  NOR2_X1 U2775 ( .A1(\mac_unit_inst/adder_reg [8]), .A2(
        \mac_unit_inst/x_mult_f_reg [8]), .ZN(n2714) );
  NOR2_X1 U2776 ( .A1(\mac_unit_inst/adder_reg [9]), .A2(
        \mac_unit_inst/x_mult_f_reg [9]), .ZN(n2715) );
  NOR2_X1 U2777 ( .A1(n2714), .A2(n2715), .ZN(n2722) );
  NOR2_X1 U2778 ( .A1(\mac_unit_inst/adder_reg [10]), .A2(
        \mac_unit_inst/x_mult_f_reg [10]), .ZN(n2726) );
  NOR2_X1 U2779 ( .A1(\mac_unit_inst/adder_reg [11]), .A2(
        \mac_unit_inst/x_mult_f_reg [11]), .ZN(n2735) );
  NOR2_X1 U2780 ( .A1(n2726), .A2(n2735), .ZN(n2626) );
  NAND2_X1 U2781 ( .A1(n2722), .A2(n2626), .ZN(n2743) );
  NAND2_X1 U2782 ( .A1(n2750), .A2(n2753), .ZN(n2629) );
  NOR2_X1 U2783 ( .A1(n2743), .A2(n2629), .ZN(n2631) );
  NAND2_X1 U2784 ( .A1(\mac_unit_inst/adder_reg [8]), .A2(
        \mac_unit_inst/x_mult_f_reg [8]), .ZN(n2713) );
  NAND2_X1 U2785 ( .A1(\mac_unit_inst/adder_reg [9]), .A2(
        \mac_unit_inst/x_mult_f_reg [9]), .ZN(n2716) );
  OAI21_X1 U2786 ( .B1(n2715), .B2(n2713), .A(n2716), .ZN(n2723) );
  NAND2_X1 U2787 ( .A1(\mac_unit_inst/adder_reg [10]), .A2(
        \mac_unit_inst/x_mult_f_reg [10]), .ZN(n2731) );
  NAND2_X1 U2788 ( .A1(\mac_unit_inst/adder_reg [11]), .A2(
        \mac_unit_inst/x_mult_f_reg [11]), .ZN(n2736) );
  OAI21_X1 U2789 ( .B1(n2735), .B2(n2731), .A(n2736), .ZN(n2625) );
  AOI21_X1 U2790 ( .B1(n2626), .B2(n2723), .A(n2625), .ZN(n2742) );
  NAND2_X1 U2791 ( .A1(\mac_unit_inst/adder_reg [12]), .A2(
        \mac_unit_inst/x_mult_f_reg [12]), .ZN(n2745) );
  INV_X1 U2792 ( .A(n2745), .ZN(n2749) );
  NAND2_X1 U2793 ( .A1(\mac_unit_inst/adder_reg [13]), .A2(
        \mac_unit_inst/x_mult_f_reg [13]), .ZN(n2752) );
  INV_X1 U2794 ( .A(n2752), .ZN(n2627) );
  AOI21_X1 U2795 ( .B1(n2753), .B2(n2749), .A(n2627), .ZN(n2628) );
  OAI21_X1 U2796 ( .B1(n2742), .B2(n2629), .A(n2628), .ZN(n2630) );
  AOI21_X1 U2797 ( .B1(n2708), .B2(n2631), .A(n2630), .ZN(n2762) );
  NOR2_X1 U2798 ( .A1(\mac_unit_inst/adder_reg [14]), .A2(
        \mac_unit_inst/x_mult_f_reg [14]), .ZN(n2758) );
  NAND2_X1 U2799 ( .A1(\mac_unit_inst/adder_reg [14]), .A2(
        \mac_unit_inst/x_mult_f_reg [14]), .ZN(n2759) );
  OAI21_X1 U2800 ( .B1(n2762), .B2(n2758), .A(n2759), .ZN(n2768) );
  OR2_X1 U2801 ( .A1(\mac_unit_inst/adder_reg [15]), .A2(
        \mac_unit_inst/x_mult_f_reg [15]), .ZN(n2766) );
  NAND2_X1 U2802 ( .A1(\mac_unit_inst/adder_reg [15]), .A2(
        \mac_unit_inst/x_mult_f_reg [15]), .ZN(n2765) );
  INV_X1 U2803 ( .A(n2765), .ZN(n2632) );
  AOI21_X1 U2804 ( .B1(n2768), .B2(n2766), .A(n2632), .ZN(n2775) );
  NOR2_X1 U2805 ( .A1(\mac_unit_inst/adder_reg [16]), .A2(
        \mac_unit_inst/x_mult_f_reg [16]), .ZN(n2771) );
  NAND2_X1 U2806 ( .A1(\mac_unit_inst/adder_reg [16]), .A2(
        \mac_unit_inst/x_mult_f_reg [16]), .ZN(n2772) );
  OAI21_X1 U2807 ( .B1(n2775), .B2(n2771), .A(n2772), .ZN(n2778) );
  FA_X1 U2808 ( .A(n3369), .B(n3325), .CI(n2633), .CO(n2634), .S(n2637) );
  NOR2_X1 U2809 ( .A1(n2637), .A2(n2634), .ZN(n2648) );
  INV_X1 U2810 ( .A(n2652), .ZN(n2636) );
  NAND2_X1 U2811 ( .A1(\ctrl_conv_output_inst/conv_start_accum ), .A2(n2815), 
        .ZN(n2635) );
  NOR2_X1 U2812 ( .A1(n2635), .A2(m_valid_y), .ZN(n2651) );
  OAI211_X1 U2813 ( .C1(n2648), .C2(n2637), .A(n2636), .B(n2651), .ZN(n2638)
         );
  OAI21_X1 U2814 ( .B1(n3369), .B2(n2785), .A(n2638), .ZN(n871) );
  INV_X1 U2815 ( .A(\ctrl_conv_output_inst/N74 ), .ZN(n3308) );
  NOR3_X1 U2816 ( .A1(n3308), .A2(conv_done), .A3(
        \ctrl_conv_output_inst/m_pre_pre_valid_y ), .ZN(n3299) );
  INV_X1 U2817 ( .A(n3299), .ZN(n3303) );
  NOR2_X1 U2818 ( .A1(n2640), .A2(n3303), .ZN(n2643) );
  OAI21_X1 U2819 ( .B1(n3331), .B2(n2639), .A(n3299), .ZN(n3305) );
  INV_X1 U2820 ( .A(n3305), .ZN(n2641) );
  NOR2_X1 U2821 ( .A1(reset), .A2(conv_done), .ZN(n2823) );
  OAI21_X1 U2822 ( .B1(n2820), .B2(n2818), .A(n2823), .ZN(n2822) );
  NOR2_X1 U2823 ( .A1(n3299), .A2(n2822), .ZN(n3300) );
  AOI21_X1 U2824 ( .B1(n2641), .B2(n2640), .A(n3300), .ZN(n3304) );
  INV_X1 U2825 ( .A(n3304), .ZN(n2642) );
  MUX2_X1 U2826 ( .A(n2643), .B(n2642), .S(fmem_addr[2]), .Z(n924) );
  NOR2_X1 U2827 ( .A1(n3331), .A2(n3305), .ZN(n2646) );
  AOI21_X1 U2828 ( .B1(n3299), .B2(n3331), .A(n3300), .ZN(n2644) );
  INV_X1 U2829 ( .A(n2644), .ZN(n2645) );
  MUX2_X1 U2830 ( .A(n2646), .B(n2645), .S(fmem_addr[1]), .Z(n925) );
  INV_X1 U2831 ( .A(n2651), .ZN(n2647) );
  NOR2_X2 U2832 ( .A1(n2648), .A2(n2647), .ZN(n2730) );
  OR2_X1 U2833 ( .A1(\mac_unit_inst/adder_reg [0]), .A2(
        \mac_unit_inst/x_mult_f_reg [0]), .ZN(n2649) );
  AND2_X1 U2834 ( .A1(n2649), .A2(n2657), .ZN(n2650) );
  NAND2_X1 U2835 ( .A1(n2730), .A2(n2650), .ZN(n2653) );
  OAI211_X1 U2836 ( .C1(n2785), .C2(n3348), .A(n2653), .B(n2783), .ZN(n890) );
  INV_X1 U2837 ( .A(n2654), .ZN(n2656) );
  NAND2_X1 U2838 ( .A1(n2656), .A2(n2655), .ZN(n2658) );
  XOR2_X1 U2839 ( .A(n2658), .B(n2657), .Z(n2659) );
  NAND2_X1 U2840 ( .A1(n2730), .A2(n2659), .ZN(n2660) );
  OAI211_X1 U2841 ( .C1(n2785), .C2(n3349), .A(n2660), .B(n2783), .ZN(n889) );
  INV_X1 U2842 ( .A(n2661), .ZN(n2668) );
  INV_X1 U2843 ( .A(n2667), .ZN(n2662) );
  NAND2_X1 U2844 ( .A1(n2662), .A2(n2666), .ZN(n2663) );
  XOR2_X1 U2845 ( .A(n2668), .B(n2663), .Z(n2664) );
  NAND2_X1 U2846 ( .A1(n2730), .A2(n2664), .ZN(n2665) );
  OAI211_X1 U2847 ( .C1(n2785), .C2(n3350), .A(n2665), .B(n2783), .ZN(n888) );
  OAI21_X1 U2848 ( .B1(n2668), .B2(n2667), .A(n2666), .ZN(n2673) );
  INV_X1 U2849 ( .A(n2669), .ZN(n2671) );
  NAND2_X1 U2850 ( .A1(n2671), .A2(n2670), .ZN(n2672) );
  XNOR2_X1 U2851 ( .A(n2673), .B(n2672), .ZN(n2674) );
  NAND2_X1 U2852 ( .A1(n2730), .A2(n2674), .ZN(n2675) );
  OAI211_X1 U2853 ( .C1(n2785), .C2(n3351), .A(n2675), .B(n2783), .ZN(n887) );
  INV_X1 U2854 ( .A(n2676), .ZN(n2693) );
  INV_X1 U2855 ( .A(n2677), .ZN(n2683) );
  NAND2_X1 U2856 ( .A1(n2683), .A2(n2681), .ZN(n2678) );
  XNOR2_X1 U2857 ( .A(n2693), .B(n2678), .ZN(n2679) );
  NAND2_X1 U2858 ( .A1(n2730), .A2(n2679), .ZN(n2680) );
  OAI211_X1 U2859 ( .C1(n2785), .C2(n3352), .A(n2680), .B(n2783), .ZN(n886) );
  INV_X1 U2860 ( .A(n2681), .ZN(n2682) );
  AOI21_X1 U2861 ( .B1(n2693), .B2(n2683), .A(n2682), .ZN(n2688) );
  INV_X1 U2862 ( .A(n2684), .ZN(n2686) );
  NAND2_X1 U2863 ( .A1(n2686), .A2(n2685), .ZN(n2687) );
  XOR2_X1 U2864 ( .A(n2688), .B(n2687), .Z(n2689) );
  NAND2_X1 U2865 ( .A1(n2730), .A2(n2689), .ZN(n2690) );
  OAI211_X1 U2866 ( .C1(n2785), .C2(n3353), .A(n2690), .B(n2783), .ZN(n885) );
  AOI21_X1 U2867 ( .B1(n2693), .B2(n2692), .A(n2691), .ZN(n2700) );
  INV_X1 U2868 ( .A(n2699), .ZN(n2694) );
  NAND2_X1 U2869 ( .A1(n2694), .A2(n2698), .ZN(n2695) );
  XOR2_X1 U2870 ( .A(n2700), .B(n2695), .Z(n2696) );
  NAND2_X1 U2871 ( .A1(n2730), .A2(n2696), .ZN(n2697) );
  OAI211_X1 U2872 ( .C1(n2785), .C2(n3354), .A(n2697), .B(n2783), .ZN(n884) );
  OAI21_X1 U2873 ( .B1(n2700), .B2(n2699), .A(n2698), .ZN(n2705) );
  INV_X1 U2874 ( .A(n2701), .ZN(n2703) );
  NAND2_X1 U2875 ( .A1(n2703), .A2(n2702), .ZN(n2704) );
  XNOR2_X1 U2876 ( .A(n2705), .B(n2704), .ZN(n2706) );
  NAND2_X1 U2877 ( .A1(n2730), .A2(n2706), .ZN(n2707) );
  OAI211_X1 U2878 ( .C1(n2785), .C2(n3355), .A(n2707), .B(n2783), .ZN(n883) );
  INV_X1 U2879 ( .A(n2708), .ZN(n2744) );
  INV_X1 U2880 ( .A(n2714), .ZN(n2709) );
  NAND2_X1 U2881 ( .A1(n2709), .A2(n2713), .ZN(n2710) );
  XOR2_X1 U2882 ( .A(n2744), .B(n2710), .Z(n2711) );
  NAND2_X1 U2883 ( .A1(n2730), .A2(n2711), .ZN(n2712) );
  OAI211_X1 U2884 ( .C1(n2785), .C2(n3356), .A(n2712), .B(n2783), .ZN(n882) );
  OAI21_X1 U2885 ( .B1(n2744), .B2(n2714), .A(n2713), .ZN(n2719) );
  INV_X1 U2886 ( .A(n2715), .ZN(n2717) );
  NAND2_X1 U2887 ( .A1(n2717), .A2(n2716), .ZN(n2718) );
  XNOR2_X1 U2888 ( .A(n2719), .B(n2718), .ZN(n2720) );
  NAND2_X1 U2889 ( .A1(n2730), .A2(n2720), .ZN(n2721) );
  OAI211_X1 U2890 ( .C1(n2785), .C2(n3357), .A(n2721), .B(n2783), .ZN(n881) );
  INV_X1 U2891 ( .A(n2722), .ZN(n2725) );
  INV_X1 U2892 ( .A(n2723), .ZN(n2724) );
  OAI21_X1 U2893 ( .B1(n2744), .B2(n2725), .A(n2724), .ZN(n2734) );
  INV_X1 U2894 ( .A(n2726), .ZN(n2733) );
  NAND2_X1 U2895 ( .A1(n2733), .A2(n2731), .ZN(n2727) );
  XNOR2_X1 U2896 ( .A(n2734), .B(n2727), .ZN(n2728) );
  NAND2_X1 U2897 ( .A1(n2730), .A2(n2728), .ZN(n2729) );
  OAI211_X1 U2898 ( .C1(n2785), .C2(n3358), .A(n2729), .B(n2783), .ZN(n880) );
  INV_X1 U2899 ( .A(n2731), .ZN(n2732) );
  AOI21_X1 U2900 ( .B1(n2734), .B2(n2733), .A(n2732), .ZN(n2739) );
  INV_X1 U2901 ( .A(n2735), .ZN(n2737) );
  NAND2_X1 U2902 ( .A1(n2737), .A2(n2736), .ZN(n2738) );
  XOR2_X1 U2903 ( .A(n2739), .B(n2738), .Z(n2740) );
  NAND2_X1 U2904 ( .A1(n2730), .A2(n2740), .ZN(n2741) );
  OAI211_X1 U2905 ( .C1(n2785), .C2(n3364), .A(n2741), .B(n2783), .ZN(n879) );
  OAI21_X1 U2906 ( .B1(n2744), .B2(n2743), .A(n2742), .ZN(n2751) );
  NAND2_X1 U2907 ( .A1(n2750), .A2(n2745), .ZN(n2746) );
  XNOR2_X1 U2908 ( .A(n2751), .B(n2746), .ZN(n2747) );
  NAND2_X1 U2909 ( .A1(n2730), .A2(n2747), .ZN(n2748) );
  OAI211_X1 U2910 ( .C1(n2785), .C2(n3359), .A(n2748), .B(n2783), .ZN(n878) );
  AOI21_X1 U2911 ( .B1(n2751), .B2(n2750), .A(n2749), .ZN(n2755) );
  NAND2_X1 U2912 ( .A1(n2753), .A2(n2752), .ZN(n2754) );
  XOR2_X1 U2913 ( .A(n2755), .B(n2754), .Z(n2756) );
  NAND2_X1 U2914 ( .A1(n2730), .A2(n2756), .ZN(n2757) );
  OAI211_X1 U2915 ( .C1(n2785), .C2(n3360), .A(n2757), .B(n2783), .ZN(n877) );
  INV_X1 U2916 ( .A(n2758), .ZN(n2760) );
  NAND2_X1 U2917 ( .A1(n2760), .A2(n2759), .ZN(n2761) );
  XOR2_X1 U2918 ( .A(n2762), .B(n2761), .Z(n2763) );
  NAND2_X1 U2919 ( .A1(n2730), .A2(n2763), .ZN(n2764) );
  OAI211_X1 U2920 ( .C1(n2785), .C2(n3361), .A(n2764), .B(n2783), .ZN(n876) );
  NAND2_X1 U2921 ( .A1(n2766), .A2(n2765), .ZN(n2767) );
  XNOR2_X1 U2922 ( .A(n2768), .B(n2767), .ZN(n2769) );
  NAND2_X1 U2923 ( .A1(n2730), .A2(n2769), .ZN(n2770) );
  OAI211_X1 U2924 ( .C1(n2785), .C2(n3362), .A(n2770), .B(n2783), .ZN(n875) );
  INV_X1 U2925 ( .A(n2771), .ZN(n2773) );
  NAND2_X1 U2926 ( .A1(n2773), .A2(n2772), .ZN(n2774) );
  XOR2_X1 U2927 ( .A(n2775), .B(n2774), .Z(n2776) );
  NAND2_X1 U2928 ( .A1(n2730), .A2(n2776), .ZN(n2777) );
  OAI211_X1 U2929 ( .C1(n2785), .C2(n3363), .A(n2777), .B(n2783), .ZN(n874) );
  FA_X1 U2930 ( .A(\mac_unit_inst/adder_reg [17]), .B(
        \mac_unit_inst/x_mult_f_reg [17]), .CI(n2778), .CO(n2781), .S(n2779)
         );
  NAND2_X1 U2931 ( .A1(n2730), .A2(n2779), .ZN(n2780) );
  OAI211_X1 U2932 ( .C1(n2785), .C2(n3365), .A(n2780), .B(n2783), .ZN(n873) );
  FA_X1 U2933 ( .A(\mac_unit_inst/adder_reg [18]), .B(
        \mac_unit_inst/x_mult_f_reg [18]), .CI(n2781), .CO(n2633), .S(n2782)
         );
  NAND2_X1 U2934 ( .A1(n2730), .A2(n2782), .ZN(n2784) );
  OAI211_X1 U2935 ( .C1(n2785), .C2(n3366), .A(n2784), .B(n2783), .ZN(n872) );
  INV_X1 U2936 ( .A(n2786), .ZN(n2787) );
  OR2_X1 U2937 ( .A1(n2788), .A2(n2787), .ZN(n2790) );
  NAND2_X1 U2938 ( .A1(n2788), .A2(n2787), .ZN(n2789) );
  NAND2_X1 U2939 ( .A1(n2790), .A2(n2789), .ZN(n2791) );
  XNOR2_X1 U2940 ( .A(n2792), .B(n2791), .ZN(n2798) );
  INV_X1 U2941 ( .A(n2794), .ZN(n2795) );
  OAI211_X1 U2942 ( .C1(n2798), .C2(n2797), .A(n2796), .B(n2795), .ZN(n2799)
         );
  OAI21_X1 U2943 ( .B1(n3325), .B2(n2800), .A(n2799), .ZN(n891) );
  NAND4_X1 U2944 ( .A1(\ctrl_conv_output_inst/cnt_conv [3]), .A2(n3333), .A3(
        n3337), .A4(n3343), .ZN(n2801) );
  NOR4_X1 U2945 ( .A1(\ctrl_conv_output_inst/cnt_conv [2]), .A2(reset), .A3(
        n2820), .A4(n2801), .ZN(\ctrl_conv_output_inst/N77 ) );
  NOR2_X1 U2947 ( .A1(s_ready_x), .A2(reset), .ZN(N29) );
  NOR2_X1 U2948 ( .A1(\ctrl_conv_output_inst/m_pre_pre_valid_y ), .A2(n2818), 
        .ZN(n2821) );
  NAND3_X1 U2949 ( .A1(n2821), .A2(n2802), .A3(n2815), .ZN(n2803) );
  OAI21_X1 U2950 ( .B1(n3307), .B2(n3344), .A(n2803), .ZN(n1339) );
  NAND2_X1 U2951 ( .A1(\ctrl_conv_output_inst/m_pre_pre_valid_y ), .A2(n3336), 
        .ZN(n2807) );
  NAND3_X1 U2952 ( .A1(\ctrl_conv_output_inst/cnt_conv [2]), .A2(
        \ctrl_conv_output_inst/cnt_conv [0]), .A3(
        \ctrl_conv_output_inst/cnt_conv [1]), .ZN(n2813) );
  OAI21_X1 U2953 ( .B1(n2807), .B2(n2813), .A(n2823), .ZN(n2814) );
  NAND3_X1 U2954 ( .A1(n3336), .A2(\ctrl_conv_output_inst/m_pre_pre_valid_y ), 
        .A3(n2823), .ZN(n2805) );
  INV_X1 U2955 ( .A(n2805), .ZN(n2808) );
  NAND2_X1 U2956 ( .A1(n2808), .A2(n3342), .ZN(n2812) );
  OR4_X1 U2957 ( .A1(n3342), .A2(n2805), .A3(n2813), .A4(
        \ctrl_conv_output_inst/cnt_conv [4]), .ZN(n2804) );
  OAI221_X1 U2958 ( .B1(n3337), .B2(n2814), .C1(n3337), .C2(n2812), .A(n2804), 
        .ZN(n1338) );
  OAI21_X1 U2959 ( .B1(\ctrl_conv_output_inst/m_pre_valid_y ), .B2(n3344), .A(
        n2823), .ZN(n2806) );
  AOI22_X1 U2960 ( .A1(\ctrl_conv_output_inst/cnt_conv [0]), .A2(n2806), .B1(
        n2805), .B2(n3333), .ZN(n1337) );
  OAI21_X1 U2961 ( .B1(n3333), .B2(n2807), .A(n2823), .ZN(n2811) );
  NAND2_X1 U2962 ( .A1(n2808), .A2(n3343), .ZN(n2810) );
  OAI22_X1 U2963 ( .A1(n2811), .A2(n3343), .B1(n3333), .B2(n2810), .ZN(n1336)
         );
  NAND4_X1 U2964 ( .A1(\ctrl_conv_output_inst/cnt_conv [0]), .A2(
        \ctrl_conv_output_inst/cnt_conv [1]), .A3(n2808), .A4(n3341), .ZN(
        n2809) );
  OAI221_X1 U2965 ( .B1(n3341), .B2(n2811), .C1(n3341), .C2(n2810), .A(n2809), 
        .ZN(n1335) );
  OAI22_X1 U2966 ( .A1(n2814), .A2(n3342), .B1(n2813), .B2(n2812), .ZN(n1334)
         );
  NAND2_X1 U2967 ( .A1(m_valid_y), .A2(n2815), .ZN(n2816) );
  OAI22_X1 U2968 ( .A1(m_ready_y), .A2(n2816), .B1(n3336), .B2(n3308), .ZN(
        n1333) );
  OAI21_X1 U2969 ( .B1(n3296), .B2(n3367), .A(n2823), .ZN(n1332) );
  NOR2_X1 U2970 ( .A1(n2820), .A2(n2818), .ZN(n2819) );
  NAND2_X1 U2971 ( .A1(n2819), .A2(n2823), .ZN(n2840) );
  AND2_X1 U2972 ( .A1(n2821), .A2(n2820), .ZN(n2824) );
  NOR3_X1 U2973 ( .A1(n2908), .A2(n2824), .A3(n2822), .ZN(n2838) );
  OAI211_X1 U2974 ( .C1(n2908), .C2(n2824), .A(n3297), .B(n2823), .ZN(n2833)
         );
  INV_X1 U2975 ( .A(n2833), .ZN(n2837) );
  AOI22_X1 U2976 ( .A1(xmem_addr[0]), .A2(n2838), .B1(n2837), .B2(n3338), .ZN(
        n2825) );
  OAI21_X1 U2977 ( .B1(n2840), .B2(n3333), .A(n2825), .ZN(n1331) );
  INV_X1 U2978 ( .A(n2840), .ZN(n2826) );
  AOI22_X1 U2979 ( .A1(n2838), .A2(xmem_addr[1]), .B1(n2826), .B2(
        \ctrl_conv_output_inst/cnt_conv [1]), .ZN(n2827) );
  OAI221_X1 U2980 ( .B1(n2833), .B2(n3137), .C1(n2833), .C2(n3160), .A(n2827), 
        .ZN(n1330) );
  XOR2_X1 U2981 ( .A(n3340), .B(n3184), .Z(n2828) );
  AOI22_X1 U2982 ( .A1(xmem_addr[2]), .A2(n2838), .B1(n2837), .B2(n2828), .ZN(
        n2829) );
  OAI21_X1 U2983 ( .B1(n2840), .B2(n3341), .A(n2829), .ZN(n1329) );
  AOI21_X1 U2984 ( .B1(n2837), .B2(n2830), .A(n2838), .ZN(n2834) );
  INV_X1 U2985 ( .A(n2831), .ZN(n2832) );
  OAI222_X1 U2986 ( .A1(n3342), .A2(n2840), .B1(n3335), .B2(n2834), .C1(n2833), 
        .C2(n2832), .ZN(n1328) );
  XOR2_X1 U2987 ( .A(xmem_addr[4]), .B(n2835), .Z(n2836) );
  AOI22_X1 U2988 ( .A1(xmem_addr[4]), .A2(n2838), .B1(n2837), .B2(n2836), .ZN(
        n2839) );
  OAI21_X1 U2989 ( .B1(n2840), .B2(n3337), .A(n2839), .ZN(n1327) );
  OAI22_X1 U2990 ( .A1(n2861), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[0][0] ), 
        .B2(n2860), .ZN(n2841) );
  INV_X1 U2991 ( .A(n2841), .ZN(n1326) );
  OAI22_X1 U2992 ( .A1(n2861), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[0][1] ), 
        .B2(n2860), .ZN(n2842) );
  INV_X1 U2993 ( .A(n2842), .ZN(n1325) );
  OAI22_X1 U2994 ( .A1(n2861), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[0][2] ), 
        .B2(n2860), .ZN(n2843) );
  INV_X1 U2995 ( .A(n2843), .ZN(n1324) );
  OAI22_X1 U2996 ( .A1(n2861), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[0][3] ), 
        .B2(n2860), .ZN(n2844) );
  INV_X1 U2997 ( .A(n2844), .ZN(n1323) );
  OAI22_X1 U2998 ( .A1(n2861), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[0][4] ), 
        .B2(n2860), .ZN(n2845) );
  INV_X1 U2999 ( .A(n2845), .ZN(n1322) );
  OAI22_X1 U3000 ( .A1(n2861), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[0][5] ), 
        .B2(n2860), .ZN(n2846) );
  INV_X1 U3001 ( .A(n2846), .ZN(n1321) );
  OAI22_X1 U3002 ( .A1(n2861), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[0][6] ), 
        .B2(n2860), .ZN(n2847) );
  INV_X1 U3003 ( .A(n2847), .ZN(n1320) );
  OAI22_X1 U3004 ( .A1(n2861), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[0][7] ), 
        .B2(n2860), .ZN(n2848) );
  INV_X1 U3005 ( .A(n2848), .ZN(n1319) );
  OAI22_X1 U3006 ( .A1(n2861), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[0][8] ), 
        .B2(n2860), .ZN(n2849) );
  INV_X1 U3007 ( .A(n2849), .ZN(n1318) );
  OAI22_X1 U3008 ( .A1(n2861), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[0][9] ), 
        .B2(n2860), .ZN(n2850) );
  INV_X1 U3009 ( .A(n2850), .ZN(n1317) );
  OAI22_X1 U3010 ( .A1(n2861), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[0][10] ), .B2(n2860), .ZN(n2851) );
  INV_X1 U3011 ( .A(n2851), .ZN(n1316) );
  OAI22_X1 U3012 ( .A1(n2861), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[0][11] ), .B2(n2860), .ZN(n2852) );
  INV_X1 U3013 ( .A(n2852), .ZN(n1315) );
  OAI22_X1 U3014 ( .A1(n2861), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[0][12] ), .B2(n2860), .ZN(n2853) );
  INV_X1 U3015 ( .A(n2853), .ZN(n1314) );
  OAI22_X1 U3016 ( .A1(n2861), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[0][13] ), .B2(n2860), .ZN(n2854) );
  INV_X1 U3017 ( .A(n2854), .ZN(n1313) );
  OAI22_X1 U3018 ( .A1(n2861), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[0][14] ), .B2(n2860), .ZN(n2855) );
  INV_X1 U3019 ( .A(n2855), .ZN(n1312) );
  OAI22_X1 U3020 ( .A1(n2861), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[0][15] ), .B2(n2860), .ZN(n2856) );
  INV_X1 U3021 ( .A(n2856), .ZN(n1311) );
  OAI22_X1 U3022 ( .A1(n2861), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[0][16] ), .B2(n2860), .ZN(n2857) );
  INV_X1 U3023 ( .A(n2857), .ZN(n1310) );
  OAI22_X1 U3024 ( .A1(n2861), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[0][17] ), .B2(n2860), .ZN(n2858) );
  INV_X1 U3025 ( .A(n2858), .ZN(n1309) );
  OAI22_X1 U3026 ( .A1(n2861), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[0][18] ), .B2(n2860), .ZN(n2859) );
  INV_X1 U3027 ( .A(n2859), .ZN(n1308) );
  OAI22_X1 U3028 ( .A1(n2861), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[0][19] ), .B2(n2860), .ZN(n2862) );
  INV_X1 U3029 ( .A(n2862), .ZN(n1307) );
  OAI22_X1 U3030 ( .A1(n2883), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[1][0] ), 
        .B2(n2882), .ZN(n2863) );
  INV_X1 U3031 ( .A(n2863), .ZN(n1306) );
  OAI22_X1 U3032 ( .A1(n2883), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[1][1] ), 
        .B2(n2882), .ZN(n2864) );
  INV_X1 U3033 ( .A(n2864), .ZN(n1305) );
  OAI22_X1 U3034 ( .A1(n2883), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[1][2] ), 
        .B2(n2882), .ZN(n2865) );
  INV_X1 U3035 ( .A(n2865), .ZN(n1304) );
  OAI22_X1 U3036 ( .A1(n2883), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[1][3] ), 
        .B2(n2882), .ZN(n2866) );
  INV_X1 U3037 ( .A(n2866), .ZN(n1303) );
  OAI22_X1 U3038 ( .A1(n2883), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[1][4] ), 
        .B2(n2882), .ZN(n2867) );
  INV_X1 U3039 ( .A(n2867), .ZN(n1302) );
  OAI22_X1 U3040 ( .A1(n2883), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[1][5] ), 
        .B2(n2882), .ZN(n2868) );
  INV_X1 U3041 ( .A(n2868), .ZN(n1301) );
  OAI22_X1 U3042 ( .A1(n2883), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[1][6] ), 
        .B2(n2882), .ZN(n2869) );
  INV_X1 U3043 ( .A(n2869), .ZN(n1300) );
  OAI22_X1 U3044 ( .A1(n2883), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[1][7] ), 
        .B2(n2882), .ZN(n2870) );
  INV_X1 U3045 ( .A(n2870), .ZN(n1299) );
  OAI22_X1 U3046 ( .A1(n2883), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[1][8] ), 
        .B2(n2882), .ZN(n2871) );
  INV_X1 U3047 ( .A(n2871), .ZN(n1298) );
  OAI22_X1 U3048 ( .A1(n2883), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[1][9] ), 
        .B2(n2882), .ZN(n2872) );
  INV_X1 U3049 ( .A(n2872), .ZN(n1297) );
  OAI22_X1 U3050 ( .A1(n2883), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[1][10] ), .B2(n2882), .ZN(n2873) );
  INV_X1 U3051 ( .A(n2873), .ZN(n1296) );
  OAI22_X1 U3052 ( .A1(n2883), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[1][11] ), .B2(n2882), .ZN(n2874) );
  INV_X1 U3053 ( .A(n2874), .ZN(n1295) );
  OAI22_X1 U3054 ( .A1(n2883), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[1][12] ), .B2(n2882), .ZN(n2875) );
  INV_X1 U3055 ( .A(n2875), .ZN(n1294) );
  OAI22_X1 U3056 ( .A1(n2883), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[1][13] ), .B2(n2882), .ZN(n2876) );
  INV_X1 U3057 ( .A(n2876), .ZN(n1293) );
  OAI22_X1 U3058 ( .A1(n2883), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[1][14] ), .B2(n2882), .ZN(n2877) );
  INV_X1 U3059 ( .A(n2877), .ZN(n1292) );
  OAI22_X1 U3060 ( .A1(n2883), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[1][15] ), .B2(n2882), .ZN(n2878) );
  INV_X1 U3061 ( .A(n2878), .ZN(n1291) );
  OAI22_X1 U3062 ( .A1(n2883), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[1][16] ), .B2(n2882), .ZN(n2879) );
  INV_X1 U3063 ( .A(n2879), .ZN(n1290) );
  OAI22_X1 U3064 ( .A1(n2883), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[1][17] ), .B2(n2882), .ZN(n2880) );
  INV_X1 U3065 ( .A(n2880), .ZN(n1289) );
  OAI22_X1 U3066 ( .A1(n2883), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[1][18] ), .B2(n2882), .ZN(n2881) );
  INV_X1 U3067 ( .A(n2881), .ZN(n1288) );
  OAI22_X1 U3068 ( .A1(n2883), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[1][19] ), .B2(n2882), .ZN(n2884) );
  INV_X1 U3069 ( .A(n2884), .ZN(n1287) );
  OAI22_X1 U3070 ( .A1(n2906), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[2][0] ), 
        .B2(n2905), .ZN(n2886) );
  INV_X1 U3071 ( .A(n2886), .ZN(n1286) );
  OAI22_X1 U3072 ( .A1(n2906), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[2][1] ), 
        .B2(n2905), .ZN(n2887) );
  INV_X1 U3073 ( .A(n2887), .ZN(n1285) );
  OAI22_X1 U3074 ( .A1(n2906), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[2][2] ), 
        .B2(n2905), .ZN(n2888) );
  INV_X1 U3075 ( .A(n2888), .ZN(n1284) );
  OAI22_X1 U3076 ( .A1(n2906), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[2][3] ), 
        .B2(n2905), .ZN(n2889) );
  INV_X1 U3077 ( .A(n2889), .ZN(n1283) );
  OAI22_X1 U3078 ( .A1(n2906), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[2][4] ), 
        .B2(n2905), .ZN(n2890) );
  INV_X1 U3079 ( .A(n2890), .ZN(n1282) );
  OAI22_X1 U3080 ( .A1(n2906), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[2][5] ), 
        .B2(n2905), .ZN(n2891) );
  INV_X1 U3081 ( .A(n2891), .ZN(n1281) );
  OAI22_X1 U3082 ( .A1(n2906), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[2][6] ), 
        .B2(n2905), .ZN(n2892) );
  INV_X1 U3083 ( .A(n2892), .ZN(n1280) );
  OAI22_X1 U3084 ( .A1(n2906), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[2][7] ), 
        .B2(n2905), .ZN(n2893) );
  INV_X1 U3085 ( .A(n2893), .ZN(n1279) );
  OAI22_X1 U3086 ( .A1(n2906), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[2][8] ), 
        .B2(n2905), .ZN(n2894) );
  INV_X1 U3087 ( .A(n2894), .ZN(n1278) );
  OAI22_X1 U3088 ( .A1(n2906), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[2][9] ), 
        .B2(n2905), .ZN(n2895) );
  INV_X1 U3089 ( .A(n2895), .ZN(n1277) );
  OAI22_X1 U3090 ( .A1(n2906), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[2][10] ), .B2(n2905), .ZN(n2896) );
  INV_X1 U3091 ( .A(n2896), .ZN(n1276) );
  OAI22_X1 U3092 ( .A1(n2906), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[2][11] ), .B2(n2905), .ZN(n2897) );
  INV_X1 U3093 ( .A(n2897), .ZN(n1275) );
  OAI22_X1 U3094 ( .A1(n2906), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[2][12] ), .B2(n2905), .ZN(n2898) );
  INV_X1 U3095 ( .A(n2898), .ZN(n1274) );
  OAI22_X1 U3096 ( .A1(n2906), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[2][13] ), .B2(n2905), .ZN(n2899) );
  INV_X1 U3097 ( .A(n2899), .ZN(n1273) );
  OAI22_X1 U3098 ( .A1(n2906), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[2][14] ), .B2(n2905), .ZN(n2900) );
  INV_X1 U3099 ( .A(n2900), .ZN(n1272) );
  OAI22_X1 U3100 ( .A1(n2906), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[2][15] ), .B2(n2905), .ZN(n2901) );
  INV_X1 U3101 ( .A(n2901), .ZN(n1271) );
  OAI22_X1 U3102 ( .A1(n2906), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[2][16] ), .B2(n2905), .ZN(n2902) );
  INV_X1 U3103 ( .A(n2902), .ZN(n1270) );
  OAI22_X1 U3104 ( .A1(n2906), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[2][17] ), .B2(n2905), .ZN(n2903) );
  INV_X1 U3105 ( .A(n2903), .ZN(n1269) );
  OAI22_X1 U3106 ( .A1(n2906), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[2][18] ), .B2(n2905), .ZN(n2904) );
  INV_X1 U3107 ( .A(n2904), .ZN(n1268) );
  OAI22_X1 U3108 ( .A1(n2906), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[2][19] ), .B2(n2905), .ZN(n2907) );
  INV_X1 U3109 ( .A(n2907), .ZN(n1267) );
  OAI22_X1 U3110 ( .A1(n2929), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[3][0] ), 
        .B2(n2928), .ZN(n2909) );
  INV_X1 U3111 ( .A(n2909), .ZN(n1266) );
  OAI22_X1 U3112 ( .A1(n2929), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[3][1] ), 
        .B2(n2928), .ZN(n2910) );
  INV_X1 U3113 ( .A(n2910), .ZN(n1265) );
  OAI22_X1 U3114 ( .A1(n2929), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[3][2] ), 
        .B2(n2928), .ZN(n2911) );
  INV_X1 U3115 ( .A(n2911), .ZN(n1264) );
  OAI22_X1 U3116 ( .A1(n2929), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[3][3] ), 
        .B2(n2928), .ZN(n2912) );
  INV_X1 U3117 ( .A(n2912), .ZN(n1263) );
  OAI22_X1 U3118 ( .A1(n2929), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[3][4] ), 
        .B2(n2928), .ZN(n2913) );
  INV_X1 U3119 ( .A(n2913), .ZN(n1262) );
  OAI22_X1 U3120 ( .A1(n2929), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[3][5] ), 
        .B2(n2928), .ZN(n2914) );
  INV_X1 U3121 ( .A(n2914), .ZN(n1261) );
  OAI22_X1 U3122 ( .A1(n2929), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[3][6] ), 
        .B2(n2928), .ZN(n2915) );
  INV_X1 U3123 ( .A(n2915), .ZN(n1260) );
  OAI22_X1 U3124 ( .A1(n2929), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[3][7] ), 
        .B2(n2928), .ZN(n2916) );
  INV_X1 U3125 ( .A(n2916), .ZN(n1259) );
  OAI22_X1 U3126 ( .A1(n2929), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[3][8] ), 
        .B2(n2928), .ZN(n2917) );
  INV_X1 U3127 ( .A(n2917), .ZN(n1258) );
  OAI22_X1 U3128 ( .A1(n2929), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[3][9] ), 
        .B2(n2928), .ZN(n2918) );
  INV_X1 U3129 ( .A(n2918), .ZN(n1257) );
  OAI22_X1 U3130 ( .A1(n2929), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[3][10] ), .B2(n2928), .ZN(n2919) );
  INV_X1 U3131 ( .A(n2919), .ZN(n1256) );
  OAI22_X1 U3132 ( .A1(n2929), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[3][11] ), .B2(n2928), .ZN(n2920) );
  INV_X1 U3133 ( .A(n2920), .ZN(n1255) );
  OAI22_X1 U3134 ( .A1(n2929), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[3][12] ), .B2(n2928), .ZN(n2921) );
  INV_X1 U3135 ( .A(n2921), .ZN(n1254) );
  OAI22_X1 U3136 ( .A1(n2929), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[3][13] ), .B2(n2928), .ZN(n2922) );
  INV_X1 U3137 ( .A(n2922), .ZN(n1253) );
  OAI22_X1 U3138 ( .A1(n2929), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[3][14] ), .B2(n2928), .ZN(n2923) );
  INV_X1 U3139 ( .A(n2923), .ZN(n1252) );
  OAI22_X1 U3140 ( .A1(n2929), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[3][15] ), .B2(n2928), .ZN(n2924) );
  INV_X1 U3141 ( .A(n2924), .ZN(n1251) );
  OAI22_X1 U3142 ( .A1(n2929), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[3][16] ), .B2(n2928), .ZN(n2925) );
  INV_X1 U3143 ( .A(n2925), .ZN(n1250) );
  OAI22_X1 U3144 ( .A1(n2929), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[3][17] ), .B2(n2928), .ZN(n2926) );
  INV_X1 U3145 ( .A(n2926), .ZN(n1249) );
  OAI22_X1 U3146 ( .A1(n2929), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[3][18] ), .B2(n2928), .ZN(n2927) );
  INV_X1 U3147 ( .A(n2927), .ZN(n1248) );
  OAI22_X1 U3148 ( .A1(n2929), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[3][19] ), .B2(n2928), .ZN(n2930) );
  INV_X1 U3149 ( .A(n2930), .ZN(n1247) );
  NOR2_X2 U3150 ( .A1(n3114), .A2(n2999), .ZN(n2952) );
  OAI22_X1 U3151 ( .A1(n2953), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[4][0] ), 
        .B2(n2952), .ZN(n2933) );
  INV_X1 U3152 ( .A(n2933), .ZN(n1246) );
  OAI22_X1 U3153 ( .A1(n2953), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[4][1] ), 
        .B2(n2952), .ZN(n2934) );
  INV_X1 U3154 ( .A(n2934), .ZN(n1245) );
  OAI22_X1 U3155 ( .A1(n2953), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[4][2] ), 
        .B2(n2952), .ZN(n2935) );
  INV_X1 U3156 ( .A(n2935), .ZN(n1244) );
  OAI22_X1 U3157 ( .A1(n2953), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[4][3] ), 
        .B2(n2952), .ZN(n2936) );
  INV_X1 U3158 ( .A(n2936), .ZN(n1243) );
  OAI22_X1 U3159 ( .A1(n2953), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[4][4] ), 
        .B2(n2952), .ZN(n2937) );
  INV_X1 U3160 ( .A(n2937), .ZN(n1242) );
  OAI22_X1 U3161 ( .A1(n2953), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[4][5] ), 
        .B2(n2952), .ZN(n2938) );
  INV_X1 U3162 ( .A(n2938), .ZN(n1241) );
  OAI22_X1 U3163 ( .A1(n2953), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[4][6] ), 
        .B2(n2952), .ZN(n2939) );
  INV_X1 U3164 ( .A(n2939), .ZN(n1240) );
  OAI22_X1 U3165 ( .A1(n2953), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[4][7] ), 
        .B2(n2952), .ZN(n2940) );
  INV_X1 U3166 ( .A(n2940), .ZN(n1239) );
  OAI22_X1 U3167 ( .A1(n2953), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[4][8] ), 
        .B2(n2952), .ZN(n2941) );
  INV_X1 U3168 ( .A(n2941), .ZN(n1238) );
  OAI22_X1 U3169 ( .A1(n2953), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[4][9] ), 
        .B2(n2952), .ZN(n2942) );
  INV_X1 U3170 ( .A(n2942), .ZN(n1237) );
  OAI22_X1 U3171 ( .A1(n2953), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[4][10] ), .B2(n2952), .ZN(n2943) );
  INV_X1 U3172 ( .A(n2943), .ZN(n1236) );
  OAI22_X1 U3173 ( .A1(n2953), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[4][11] ), .B2(n2952), .ZN(n2944) );
  INV_X1 U3174 ( .A(n2944), .ZN(n1235) );
  OAI22_X1 U3175 ( .A1(n2953), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[4][12] ), .B2(n2952), .ZN(n2945) );
  INV_X1 U3176 ( .A(n2945), .ZN(n1234) );
  OAI22_X1 U3177 ( .A1(n2953), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[4][13] ), .B2(n2952), .ZN(n2946) );
  INV_X1 U3178 ( .A(n2946), .ZN(n1233) );
  OAI22_X1 U3179 ( .A1(n2953), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[4][14] ), .B2(n2952), .ZN(n2947) );
  INV_X1 U3180 ( .A(n2947), .ZN(n1232) );
  OAI22_X1 U3181 ( .A1(n2953), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[4][15] ), .B2(n2952), .ZN(n2948) );
  INV_X1 U3182 ( .A(n2948), .ZN(n1231) );
  OAI22_X1 U3183 ( .A1(n2953), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[4][16] ), .B2(n2952), .ZN(n2949) );
  INV_X1 U3184 ( .A(n2949), .ZN(n1230) );
  OAI22_X1 U3185 ( .A1(n2953), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[4][17] ), .B2(n2952), .ZN(n2950) );
  INV_X1 U3186 ( .A(n2950), .ZN(n1229) );
  OAI22_X1 U3187 ( .A1(n2953), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[4][18] ), .B2(n2952), .ZN(n2951) );
  INV_X1 U3188 ( .A(n2951), .ZN(n1228) );
  OAI22_X1 U3189 ( .A1(n2953), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[4][19] ), .B2(n2952), .ZN(n2954) );
  INV_X1 U3190 ( .A(n2954), .ZN(n1227) );
  NOR2_X2 U3191 ( .A1(n3137), .A2(n2999), .ZN(n2974) );
  OAI22_X1 U3192 ( .A1(n2975), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[5][0] ), 
        .B2(n2974), .ZN(n2955) );
  INV_X1 U3193 ( .A(n2955), .ZN(n1226) );
  OAI22_X1 U3194 ( .A1(n2975), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[5][1] ), 
        .B2(n2974), .ZN(n2956) );
  INV_X1 U3195 ( .A(n2956), .ZN(n1225) );
  OAI22_X1 U3196 ( .A1(n2975), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[5][2] ), 
        .B2(n2974), .ZN(n2957) );
  INV_X1 U3197 ( .A(n2957), .ZN(n1224) );
  OAI22_X1 U3198 ( .A1(n2975), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[5][3] ), 
        .B2(n2974), .ZN(n2958) );
  INV_X1 U3199 ( .A(n2958), .ZN(n1223) );
  OAI22_X1 U3200 ( .A1(n2975), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[5][4] ), 
        .B2(n2974), .ZN(n2959) );
  INV_X1 U3201 ( .A(n2959), .ZN(n1222) );
  OAI22_X1 U3202 ( .A1(n2975), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[5][5] ), 
        .B2(n2974), .ZN(n2960) );
  INV_X1 U3203 ( .A(n2960), .ZN(n1221) );
  OAI22_X1 U3204 ( .A1(n2975), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[5][6] ), 
        .B2(n2974), .ZN(n2961) );
  INV_X1 U3205 ( .A(n2961), .ZN(n1220) );
  OAI22_X1 U3206 ( .A1(n2975), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[5][7] ), 
        .B2(n2974), .ZN(n2962) );
  INV_X1 U3207 ( .A(n2962), .ZN(n1219) );
  OAI22_X1 U3208 ( .A1(n2975), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[5][8] ), 
        .B2(n2974), .ZN(n2963) );
  INV_X1 U3209 ( .A(n2963), .ZN(n1218) );
  OAI22_X1 U3210 ( .A1(n2975), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[5][9] ), 
        .B2(n2974), .ZN(n2964) );
  INV_X1 U3211 ( .A(n2964), .ZN(n1217) );
  OAI22_X1 U3212 ( .A1(n2975), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[5][10] ), .B2(n2974), .ZN(n2965) );
  INV_X1 U3213 ( .A(n2965), .ZN(n1216) );
  OAI22_X1 U3214 ( .A1(n2975), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[5][11] ), .B2(n2974), .ZN(n2966) );
  INV_X1 U3215 ( .A(n2966), .ZN(n1215) );
  OAI22_X1 U3216 ( .A1(n2975), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[5][12] ), .B2(n2974), .ZN(n2967) );
  INV_X1 U3217 ( .A(n2967), .ZN(n1214) );
  OAI22_X1 U3218 ( .A1(n2975), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[5][13] ), .B2(n2974), .ZN(n2968) );
  INV_X1 U3219 ( .A(n2968), .ZN(n1213) );
  OAI22_X1 U3220 ( .A1(n2975), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[5][14] ), .B2(n2974), .ZN(n2969) );
  INV_X1 U3221 ( .A(n2969), .ZN(n1212) );
  OAI22_X1 U3222 ( .A1(n2975), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[5][15] ), .B2(n2974), .ZN(n2970) );
  INV_X1 U3223 ( .A(n2970), .ZN(n1211) );
  OAI22_X1 U3224 ( .A1(n2975), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[5][16] ), .B2(n2974), .ZN(n2971) );
  INV_X1 U3225 ( .A(n2971), .ZN(n1210) );
  OAI22_X1 U3226 ( .A1(n2975), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[5][17] ), .B2(n2974), .ZN(n2972) );
  INV_X1 U3227 ( .A(n2972), .ZN(n1209) );
  OAI22_X1 U3228 ( .A1(n2975), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[5][18] ), .B2(n2974), .ZN(n2973) );
  INV_X1 U3229 ( .A(n2973), .ZN(n1208) );
  OAI22_X1 U3230 ( .A1(n2975), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[5][19] ), .B2(n2974), .ZN(n2976) );
  INV_X1 U3231 ( .A(n2976), .ZN(n1207) );
  NOR2_X2 U3232 ( .A1(n3160), .A2(n2999), .ZN(n2996) );
  OAI22_X1 U3233 ( .A1(n2997), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[6][0] ), 
        .B2(n2996), .ZN(n2977) );
  INV_X1 U3234 ( .A(n2977), .ZN(n1206) );
  OAI22_X1 U3235 ( .A1(n2997), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[6][1] ), 
        .B2(n2996), .ZN(n2978) );
  INV_X1 U3236 ( .A(n2978), .ZN(n1205) );
  OAI22_X1 U3237 ( .A1(n2997), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[6][2] ), 
        .B2(n2996), .ZN(n2979) );
  INV_X1 U3238 ( .A(n2979), .ZN(n1204) );
  OAI22_X1 U3239 ( .A1(n2997), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[6][3] ), 
        .B2(n2996), .ZN(n2980) );
  INV_X1 U3240 ( .A(n2980), .ZN(n1203) );
  OAI22_X1 U3241 ( .A1(n2997), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[6][4] ), 
        .B2(n2996), .ZN(n2981) );
  INV_X1 U3242 ( .A(n2981), .ZN(n1202) );
  OAI22_X1 U3243 ( .A1(n2997), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[6][5] ), 
        .B2(n2996), .ZN(n2982) );
  INV_X1 U3244 ( .A(n2982), .ZN(n1201) );
  OAI22_X1 U3245 ( .A1(n2997), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[6][6] ), 
        .B2(n2996), .ZN(n2983) );
  INV_X1 U3246 ( .A(n2983), .ZN(n1200) );
  OAI22_X1 U3247 ( .A1(n2997), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[6][7] ), 
        .B2(n2996), .ZN(n2984) );
  INV_X1 U3248 ( .A(n2984), .ZN(n1199) );
  OAI22_X1 U3249 ( .A1(n2997), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[6][8] ), 
        .B2(n2996), .ZN(n2985) );
  INV_X1 U3250 ( .A(n2985), .ZN(n1198) );
  OAI22_X1 U3251 ( .A1(n2997), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[6][9] ), 
        .B2(n2996), .ZN(n2986) );
  INV_X1 U3252 ( .A(n2986), .ZN(n1197) );
  OAI22_X1 U3253 ( .A1(n2997), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[6][10] ), .B2(n2996), .ZN(n2987) );
  INV_X1 U3254 ( .A(n2987), .ZN(n1196) );
  OAI22_X1 U3255 ( .A1(n2997), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[6][11] ), .B2(n2996), .ZN(n2988) );
  INV_X1 U3256 ( .A(n2988), .ZN(n1195) );
  OAI22_X1 U3257 ( .A1(n2997), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[6][12] ), .B2(n2996), .ZN(n2989) );
  INV_X1 U3258 ( .A(n2989), .ZN(n1194) );
  OAI22_X1 U3259 ( .A1(n2997), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[6][13] ), .B2(n2996), .ZN(n2990) );
  INV_X1 U3260 ( .A(n2990), .ZN(n1193) );
  OAI22_X1 U3261 ( .A1(n2997), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[6][14] ), .B2(n2996), .ZN(n2991) );
  INV_X1 U3262 ( .A(n2991), .ZN(n1192) );
  OAI22_X1 U3263 ( .A1(n2997), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[6][15] ), .B2(n2996), .ZN(n2992) );
  INV_X1 U3264 ( .A(n2992), .ZN(n1191) );
  OAI22_X1 U3265 ( .A1(n2997), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[6][16] ), .B2(n2996), .ZN(n2993) );
  INV_X1 U3266 ( .A(n2993), .ZN(n1190) );
  OAI22_X1 U3267 ( .A1(n2997), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[6][17] ), .B2(n2996), .ZN(n2994) );
  INV_X1 U3268 ( .A(n2994), .ZN(n1189) );
  OAI22_X1 U3269 ( .A1(n2997), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[6][18] ), .B2(n2996), .ZN(n2995) );
  INV_X1 U3270 ( .A(n2995), .ZN(n1188) );
  OAI22_X1 U3271 ( .A1(n2997), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[6][19] ), .B2(n2996), .ZN(n2998) );
  INV_X1 U3272 ( .A(n2998), .ZN(n1187) );
  NOR2_X2 U3273 ( .A1(n3184), .A2(n2999), .ZN(n3019) );
  OAI22_X1 U3274 ( .A1(n3020), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[7][0] ), 
        .B2(n3019), .ZN(n3000) );
  INV_X1 U3275 ( .A(n3000), .ZN(n1186) );
  OAI22_X1 U3276 ( .A1(n3020), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[7][1] ), 
        .B2(n3019), .ZN(n3001) );
  INV_X1 U3277 ( .A(n3001), .ZN(n1185) );
  OAI22_X1 U3278 ( .A1(n3020), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[7][2] ), 
        .B2(n3019), .ZN(n3002) );
  INV_X1 U3279 ( .A(n3002), .ZN(n1184) );
  OAI22_X1 U3280 ( .A1(n3020), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[7][3] ), 
        .B2(n3019), .ZN(n3003) );
  INV_X1 U3281 ( .A(n3003), .ZN(n1183) );
  OAI22_X1 U3282 ( .A1(n3020), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[7][4] ), 
        .B2(n3019), .ZN(n3004) );
  INV_X1 U3283 ( .A(n3004), .ZN(n1182) );
  OAI22_X1 U3284 ( .A1(n3020), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[7][5] ), 
        .B2(n3019), .ZN(n3005) );
  INV_X1 U3285 ( .A(n3005), .ZN(n1181) );
  OAI22_X1 U3286 ( .A1(n3020), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[7][6] ), 
        .B2(n3019), .ZN(n3006) );
  INV_X1 U3287 ( .A(n3006), .ZN(n1180) );
  OAI22_X1 U3288 ( .A1(n3020), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[7][7] ), 
        .B2(n3019), .ZN(n3007) );
  INV_X1 U3289 ( .A(n3007), .ZN(n1179) );
  OAI22_X1 U3290 ( .A1(n3020), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[7][8] ), 
        .B2(n3019), .ZN(n3008) );
  INV_X1 U3291 ( .A(n3008), .ZN(n1178) );
  OAI22_X1 U3292 ( .A1(n3020), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[7][9] ), 
        .B2(n3019), .ZN(n3009) );
  INV_X1 U3293 ( .A(n3009), .ZN(n1177) );
  OAI22_X1 U3294 ( .A1(n3020), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[7][10] ), .B2(n3019), .ZN(n3010) );
  INV_X1 U3295 ( .A(n3010), .ZN(n1176) );
  OAI22_X1 U3296 ( .A1(n3020), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[7][11] ), .B2(n3019), .ZN(n3011) );
  INV_X1 U3297 ( .A(n3011), .ZN(n1175) );
  OAI22_X1 U3298 ( .A1(n3020), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[7][12] ), .B2(n3019), .ZN(n3012) );
  INV_X1 U3299 ( .A(n3012), .ZN(n1174) );
  OAI22_X1 U3300 ( .A1(n3020), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[7][13] ), .B2(n3019), .ZN(n3013) );
  INV_X1 U3301 ( .A(n3013), .ZN(n1173) );
  OAI22_X1 U3302 ( .A1(n3020), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[7][14] ), .B2(n3019), .ZN(n3014) );
  INV_X1 U3303 ( .A(n3014), .ZN(n1172) );
  OAI22_X1 U3304 ( .A1(n3020), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[7][15] ), .B2(n3019), .ZN(n3015) );
  INV_X1 U3305 ( .A(n3015), .ZN(n1171) );
  OAI22_X1 U3306 ( .A1(n3020), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[7][16] ), .B2(n3019), .ZN(n3016) );
  INV_X1 U3307 ( .A(n3016), .ZN(n1170) );
  OAI22_X1 U3308 ( .A1(n3020), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[7][17] ), .B2(n3019), .ZN(n3017) );
  INV_X1 U3309 ( .A(n3017), .ZN(n1169) );
  OAI22_X1 U3310 ( .A1(n3020), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[7][18] ), .B2(n3019), .ZN(n3018) );
  INV_X1 U3311 ( .A(n3018), .ZN(n1168) );
  OAI22_X1 U3312 ( .A1(n3020), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[7][19] ), .B2(n3019), .ZN(n3021) );
  INV_X1 U3313 ( .A(n3021), .ZN(n1167) );
  NAND2_X1 U3314 ( .A1(n3022), .A2(n3112), .ZN(n3089) );
  OAI22_X1 U3315 ( .A1(n3043), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[8][0] ), 
        .B2(n3042), .ZN(n3023) );
  INV_X1 U3316 ( .A(n3023), .ZN(n1166) );
  OAI22_X1 U3317 ( .A1(n3043), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[8][1] ), 
        .B2(n3042), .ZN(n3024) );
  INV_X1 U3318 ( .A(n3024), .ZN(n1165) );
  OAI22_X1 U3319 ( .A1(n3043), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[8][2] ), 
        .B2(n3042), .ZN(n3025) );
  INV_X1 U3320 ( .A(n3025), .ZN(n1164) );
  OAI22_X1 U3321 ( .A1(n3043), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[8][3] ), 
        .B2(n3042), .ZN(n3026) );
  INV_X1 U3322 ( .A(n3026), .ZN(n1163) );
  OAI22_X1 U3323 ( .A1(n3043), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[8][4] ), 
        .B2(n3042), .ZN(n3027) );
  INV_X1 U3324 ( .A(n3027), .ZN(n1162) );
  OAI22_X1 U3325 ( .A1(n3043), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[8][5] ), 
        .B2(n3042), .ZN(n3028) );
  INV_X1 U3326 ( .A(n3028), .ZN(n1161) );
  OAI22_X1 U3327 ( .A1(n3043), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[8][6] ), 
        .B2(n3042), .ZN(n3029) );
  INV_X1 U3328 ( .A(n3029), .ZN(n1160) );
  OAI22_X1 U3329 ( .A1(n3043), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[8][7] ), 
        .B2(n3042), .ZN(n3030) );
  INV_X1 U3330 ( .A(n3030), .ZN(n1159) );
  OAI22_X1 U3331 ( .A1(n3043), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[8][8] ), 
        .B2(n3042), .ZN(n3031) );
  INV_X1 U3332 ( .A(n3031), .ZN(n1158) );
  OAI22_X1 U3333 ( .A1(n3043), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[8][9] ), 
        .B2(n3042), .ZN(n3032) );
  INV_X1 U3334 ( .A(n3032), .ZN(n1157) );
  OAI22_X1 U3335 ( .A1(n3043), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[8][10] ), .B2(n3042), .ZN(n3033) );
  INV_X1 U3336 ( .A(n3033), .ZN(n1156) );
  OAI22_X1 U3337 ( .A1(n3043), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[8][11] ), .B2(n3042), .ZN(n3034) );
  INV_X1 U3338 ( .A(n3034), .ZN(n1155) );
  OAI22_X1 U3339 ( .A1(n3043), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[8][12] ), .B2(n3042), .ZN(n3035) );
  INV_X1 U3340 ( .A(n3035), .ZN(n1154) );
  OAI22_X1 U3341 ( .A1(n3043), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[8][13] ), .B2(n3042), .ZN(n3036) );
  INV_X1 U3342 ( .A(n3036), .ZN(n1153) );
  OAI22_X1 U3343 ( .A1(n3043), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[8][14] ), .B2(n3042), .ZN(n3037) );
  INV_X1 U3344 ( .A(n3037), .ZN(n1152) );
  OAI22_X1 U3345 ( .A1(n3043), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[8][15] ), .B2(n3042), .ZN(n3038) );
  INV_X1 U3346 ( .A(n3038), .ZN(n1151) );
  OAI22_X1 U3347 ( .A1(n3043), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[8][16] ), .B2(n3042), .ZN(n3039) );
  INV_X1 U3348 ( .A(n3039), .ZN(n1150) );
  OAI22_X1 U3349 ( .A1(n3043), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[8][17] ), .B2(n3042), .ZN(n3040) );
  INV_X1 U3350 ( .A(n3040), .ZN(n1149) );
  OAI22_X1 U3351 ( .A1(n3043), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[8][18] ), .B2(n3042), .ZN(n3041) );
  INV_X1 U3352 ( .A(n3041), .ZN(n1148) );
  OAI22_X1 U3353 ( .A1(n3043), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[8][19] ), .B2(n3042), .ZN(n3044) );
  INV_X1 U3354 ( .A(n3044), .ZN(n1147) );
  OAI22_X1 U3355 ( .A1(n3065), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[9][0] ), 
        .B2(n3045), .ZN(n3046) );
  INV_X1 U3356 ( .A(n3046), .ZN(n1146) );
  OAI22_X1 U3357 ( .A1(n3065), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[9][1] ), 
        .B2(n3045), .ZN(n3047) );
  INV_X1 U3358 ( .A(n3047), .ZN(n1145) );
  OAI22_X1 U3359 ( .A1(n3065), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[9][2] ), 
        .B2(n3045), .ZN(n3048) );
  INV_X1 U3360 ( .A(n3048), .ZN(n1144) );
  OAI22_X1 U3361 ( .A1(n3065), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[9][3] ), 
        .B2(n3045), .ZN(n3049) );
  INV_X1 U3362 ( .A(n3049), .ZN(n1143) );
  OAI22_X1 U3363 ( .A1(n3065), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[9][4] ), 
        .B2(n3045), .ZN(n3050) );
  INV_X1 U3364 ( .A(n3050), .ZN(n1142) );
  OAI22_X1 U3365 ( .A1(n3065), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[9][5] ), 
        .B2(n3045), .ZN(n3051) );
  INV_X1 U3366 ( .A(n3051), .ZN(n1141) );
  OAI22_X1 U3367 ( .A1(n3065), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[9][6] ), 
        .B2(n3045), .ZN(n3052) );
  INV_X1 U3368 ( .A(n3052), .ZN(n1140) );
  OAI22_X1 U3369 ( .A1(n3065), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[9][7] ), 
        .B2(n3045), .ZN(n3053) );
  INV_X1 U3370 ( .A(n3053), .ZN(n1139) );
  OAI22_X1 U3371 ( .A1(n3065), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[9][8] ), 
        .B2(n3045), .ZN(n3054) );
  INV_X1 U3372 ( .A(n3054), .ZN(n1138) );
  OAI22_X1 U3373 ( .A1(n3065), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[9][9] ), 
        .B2(n3045), .ZN(n3055) );
  INV_X1 U3374 ( .A(n3055), .ZN(n1137) );
  OAI22_X1 U3375 ( .A1(n3065), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[9][10] ), .B2(n3045), .ZN(n3056) );
  INV_X1 U3376 ( .A(n3056), .ZN(n1136) );
  OAI22_X1 U3377 ( .A1(n3065), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[9][11] ), .B2(n3045), .ZN(n3057) );
  INV_X1 U3378 ( .A(n3057), .ZN(n1135) );
  OAI22_X1 U3379 ( .A1(n3065), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[9][12] ), .B2(n3045), .ZN(n3058) );
  INV_X1 U3380 ( .A(n3058), .ZN(n1134) );
  OAI22_X1 U3381 ( .A1(n3065), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[9][13] ), .B2(n3045), .ZN(n3059) );
  INV_X1 U3382 ( .A(n3059), .ZN(n1133) );
  OAI22_X1 U3383 ( .A1(n3065), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[9][14] ), .B2(n3045), .ZN(n3060) );
  INV_X1 U3384 ( .A(n3060), .ZN(n1132) );
  OAI22_X1 U3385 ( .A1(n3065), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[9][15] ), .B2(n3045), .ZN(n3061) );
  INV_X1 U3386 ( .A(n3061), .ZN(n1131) );
  OAI22_X1 U3387 ( .A1(n3065), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[9][16] ), .B2(n3045), .ZN(n3062) );
  INV_X1 U3388 ( .A(n3062), .ZN(n1130) );
  OAI22_X1 U3389 ( .A1(n3065), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[9][17] ), .B2(n3045), .ZN(n3063) );
  INV_X1 U3390 ( .A(n3063), .ZN(n1129) );
  OAI22_X1 U3391 ( .A1(n3065), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[9][18] ), .B2(n3045), .ZN(n3064) );
  INV_X1 U3392 ( .A(n3064), .ZN(n1128) );
  OAI22_X1 U3393 ( .A1(n3065), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[9][19] ), .B2(n3045), .ZN(n3066) );
  INV_X1 U3394 ( .A(n3066), .ZN(n1127) );
  OAI22_X1 U3395 ( .A1(n3087), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[10][0] ), .B2(n3067), .ZN(n3068) );
  INV_X1 U3396 ( .A(n3068), .ZN(n1126) );
  OAI22_X1 U3397 ( .A1(n3087), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[10][1] ), .B2(n3067), .ZN(n3069) );
  INV_X1 U3398 ( .A(n3069), .ZN(n1125) );
  OAI22_X1 U3399 ( .A1(n3087), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[10][2] ), .B2(n3067), .ZN(n3070) );
  INV_X1 U3400 ( .A(n3070), .ZN(n1124) );
  OAI22_X1 U3401 ( .A1(n3087), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[10][3] ), .B2(n3067), .ZN(n3071) );
  INV_X1 U3402 ( .A(n3071), .ZN(n1123) );
  OAI22_X1 U3403 ( .A1(n3087), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[10][4] ), .B2(n3067), .ZN(n3072) );
  INV_X1 U3404 ( .A(n3072), .ZN(n1122) );
  OAI22_X1 U3405 ( .A1(n3087), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[10][5] ), .B2(n3067), .ZN(n3073) );
  INV_X1 U3406 ( .A(n3073), .ZN(n1121) );
  OAI22_X1 U3407 ( .A1(n3087), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[10][6] ), .B2(n3067), .ZN(n3074) );
  INV_X1 U3408 ( .A(n3074), .ZN(n1120) );
  OAI22_X1 U3409 ( .A1(n3087), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[10][7] ), .B2(n3067), .ZN(n3075) );
  INV_X1 U3410 ( .A(n3075), .ZN(n1119) );
  OAI22_X1 U3411 ( .A1(n3087), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[10][8] ), .B2(n3067), .ZN(n3076) );
  INV_X1 U3412 ( .A(n3076), .ZN(n1118) );
  OAI22_X1 U3413 ( .A1(n3087), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[10][9] ), .B2(n3067), .ZN(n3077) );
  INV_X1 U3414 ( .A(n3077), .ZN(n1117) );
  OAI22_X1 U3415 ( .A1(n3087), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[10][10] ), .B2(n3067), .ZN(n3078) );
  INV_X1 U3416 ( .A(n3078), .ZN(n1116) );
  OAI22_X1 U3417 ( .A1(n3087), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[10][11] ), .B2(n3067), .ZN(n3079) );
  INV_X1 U3418 ( .A(n3079), .ZN(n1115) );
  OAI22_X1 U3419 ( .A1(n3087), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[10][12] ), .B2(n3067), .ZN(n3080) );
  INV_X1 U3420 ( .A(n3080), .ZN(n1114) );
  OAI22_X1 U3421 ( .A1(n3087), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[10][13] ), .B2(n3067), .ZN(n3081) );
  INV_X1 U3422 ( .A(n3081), .ZN(n1113) );
  OAI22_X1 U3423 ( .A1(n3087), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[10][14] ), .B2(n3067), .ZN(n3082) );
  INV_X1 U3424 ( .A(n3082), .ZN(n1112) );
  OAI22_X1 U3425 ( .A1(n3087), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[10][15] ), .B2(n3067), .ZN(n3083) );
  INV_X1 U3426 ( .A(n3083), .ZN(n1111) );
  OAI22_X1 U3427 ( .A1(n3087), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[10][16] ), .B2(n3067), .ZN(n3084) );
  INV_X1 U3428 ( .A(n3084), .ZN(n1110) );
  OAI22_X1 U3429 ( .A1(n3087), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[10][17] ), .B2(n3067), .ZN(n3085) );
  INV_X1 U3430 ( .A(n3085), .ZN(n1109) );
  OAI22_X1 U3431 ( .A1(n3087), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[10][18] ), .B2(n3067), .ZN(n3086) );
  INV_X1 U3432 ( .A(n3086), .ZN(n1108) );
  OAI22_X1 U3433 ( .A1(n3087), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[10][19] ), .B2(n3067), .ZN(n3088) );
  INV_X1 U3434 ( .A(n3088), .ZN(n1107) );
  OAI22_X1 U3435 ( .A1(n3110), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[11][0] ), .B2(n3090), .ZN(n3091) );
  INV_X1 U3436 ( .A(n3091), .ZN(n1106) );
  OAI22_X1 U3437 ( .A1(n3110), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[11][1] ), .B2(n3090), .ZN(n3092) );
  INV_X1 U3438 ( .A(n3092), .ZN(n1105) );
  OAI22_X1 U3439 ( .A1(n3110), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[11][2] ), .B2(n3090), .ZN(n3093) );
  INV_X1 U3440 ( .A(n3093), .ZN(n1104) );
  OAI22_X1 U3441 ( .A1(n3110), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[11][3] ), .B2(n3090), .ZN(n3094) );
  INV_X1 U3442 ( .A(n3094), .ZN(n1103) );
  OAI22_X1 U3443 ( .A1(n3110), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[11][4] ), .B2(n3090), .ZN(n3095) );
  INV_X1 U3444 ( .A(n3095), .ZN(n1102) );
  OAI22_X1 U3445 ( .A1(n3110), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[11][5] ), .B2(n3090), .ZN(n3096) );
  INV_X1 U3446 ( .A(n3096), .ZN(n1101) );
  OAI22_X1 U3447 ( .A1(n3110), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[11][6] ), .B2(n3090), .ZN(n3097) );
  INV_X1 U3448 ( .A(n3097), .ZN(n1100) );
  OAI22_X1 U3449 ( .A1(n3110), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[11][7] ), .B2(n3090), .ZN(n3098) );
  INV_X1 U3450 ( .A(n3098), .ZN(n1099) );
  OAI22_X1 U3451 ( .A1(n3110), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[11][8] ), .B2(n3090), .ZN(n3099) );
  INV_X1 U3452 ( .A(n3099), .ZN(n1098) );
  OAI22_X1 U3453 ( .A1(n3110), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[11][9] ), .B2(n3090), .ZN(n3100) );
  INV_X1 U3454 ( .A(n3100), .ZN(n1097) );
  OAI22_X1 U3455 ( .A1(n3110), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[11][10] ), .B2(n3090), .ZN(n3101) );
  INV_X1 U3456 ( .A(n3101), .ZN(n1096) );
  OAI22_X1 U3457 ( .A1(n3110), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[11][11] ), .B2(n3090), .ZN(n3102) );
  INV_X1 U3458 ( .A(n3102), .ZN(n1095) );
  OAI22_X1 U3459 ( .A1(n3110), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[11][12] ), .B2(n3090), .ZN(n3103) );
  INV_X1 U3460 ( .A(n3103), .ZN(n1094) );
  OAI22_X1 U3461 ( .A1(n3110), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[11][13] ), .B2(n3090), .ZN(n3104) );
  INV_X1 U3462 ( .A(n3104), .ZN(n1093) );
  OAI22_X1 U3463 ( .A1(n3110), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[11][14] ), .B2(n3090), .ZN(n3105) );
  INV_X1 U3464 ( .A(n3105), .ZN(n1092) );
  OAI22_X1 U3465 ( .A1(n3110), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[11][15] ), .B2(n3090), .ZN(n3106) );
  INV_X1 U3466 ( .A(n3106), .ZN(n1091) );
  OAI22_X1 U3467 ( .A1(n3110), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[11][16] ), .B2(n3090), .ZN(n3107) );
  INV_X1 U3468 ( .A(n3107), .ZN(n1090) );
  OAI22_X1 U3469 ( .A1(n3110), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[11][17] ), .B2(n3090), .ZN(n3108) );
  INV_X1 U3470 ( .A(n3108), .ZN(n1089) );
  OAI22_X1 U3471 ( .A1(n3110), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[11][18] ), .B2(n3090), .ZN(n3109) );
  INV_X1 U3472 ( .A(n3109), .ZN(n1088) );
  OAI22_X1 U3473 ( .A1(n3110), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[11][19] ), .B2(n3090), .ZN(n3111) );
  INV_X1 U3474 ( .A(n3111), .ZN(n1087) );
  NAND2_X1 U3475 ( .A1(n3113), .A2(n3112), .ZN(n3183) );
  NOR2_X2 U3476 ( .A1(n3114), .A2(n3183), .ZN(n3134) );
  OAI22_X1 U3477 ( .A1(n3135), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[12][0] ), .B2(n3134), .ZN(n3115) );
  INV_X1 U3478 ( .A(n3115), .ZN(n1086) );
  OAI22_X1 U3479 ( .A1(n3135), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[12][1] ), .B2(n3134), .ZN(n3116) );
  INV_X1 U3480 ( .A(n3116), .ZN(n1085) );
  OAI22_X1 U3481 ( .A1(n3135), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[12][2] ), .B2(n3134), .ZN(n3117) );
  INV_X1 U3482 ( .A(n3117), .ZN(n1084) );
  OAI22_X1 U3483 ( .A1(n3135), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[12][3] ), .B2(n3134), .ZN(n3118) );
  INV_X1 U3484 ( .A(n3118), .ZN(n1083) );
  OAI22_X1 U3485 ( .A1(n3135), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[12][4] ), .B2(n3134), .ZN(n3119) );
  INV_X1 U3486 ( .A(n3119), .ZN(n1082) );
  OAI22_X1 U3487 ( .A1(n3135), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[12][5] ), .B2(n3134), .ZN(n3120) );
  INV_X1 U3488 ( .A(n3120), .ZN(n1081) );
  OAI22_X1 U3489 ( .A1(n3135), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[12][6] ), .B2(n3134), .ZN(n3121) );
  INV_X1 U3490 ( .A(n3121), .ZN(n1080) );
  OAI22_X1 U3491 ( .A1(n3135), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[12][7] ), .B2(n3134), .ZN(n3122) );
  INV_X1 U3492 ( .A(n3122), .ZN(n1079) );
  OAI22_X1 U3493 ( .A1(n3135), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[12][8] ), .B2(n3134), .ZN(n3123) );
  INV_X1 U3494 ( .A(n3123), .ZN(n1078) );
  OAI22_X1 U3495 ( .A1(n3135), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[12][9] ), .B2(n3134), .ZN(n3124) );
  INV_X1 U3496 ( .A(n3124), .ZN(n1077) );
  OAI22_X1 U3497 ( .A1(n3135), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[12][10] ), .B2(n3134), .ZN(n3125) );
  INV_X1 U3498 ( .A(n3125), .ZN(n1076) );
  OAI22_X1 U3499 ( .A1(n3135), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[12][11] ), .B2(n3134), .ZN(n3126) );
  INV_X1 U3500 ( .A(n3126), .ZN(n1075) );
  OAI22_X1 U3501 ( .A1(n3135), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[12][12] ), .B2(n3134), .ZN(n3127) );
  INV_X1 U3502 ( .A(n3127), .ZN(n1074) );
  OAI22_X1 U3503 ( .A1(n3135), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[12][13] ), .B2(n3134), .ZN(n3128) );
  INV_X1 U3504 ( .A(n3128), .ZN(n1073) );
  OAI22_X1 U3505 ( .A1(n3135), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[12][14] ), .B2(n3134), .ZN(n3129) );
  INV_X1 U3506 ( .A(n3129), .ZN(n1072) );
  OAI22_X1 U3507 ( .A1(n3135), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[12][15] ), .B2(n3134), .ZN(n3130) );
  INV_X1 U3508 ( .A(n3130), .ZN(n1071) );
  OAI22_X1 U3509 ( .A1(n3135), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[12][16] ), .B2(n3134), .ZN(n3131) );
  INV_X1 U3510 ( .A(n3131), .ZN(n1070) );
  OAI22_X1 U3511 ( .A1(n3135), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[12][17] ), .B2(n3134), .ZN(n3132) );
  INV_X1 U3512 ( .A(n3132), .ZN(n1069) );
  OAI22_X1 U3513 ( .A1(n3135), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[12][18] ), .B2(n3134), .ZN(n3133) );
  INV_X1 U3514 ( .A(n3133), .ZN(n1068) );
  OAI22_X1 U3515 ( .A1(n3135), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[12][19] ), .B2(n3134), .ZN(n3136) );
  INV_X1 U3516 ( .A(n3136), .ZN(n1067) );
  OAI22_X1 U3517 ( .A1(n3158), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[13][0] ), .B2(n3157), .ZN(n3138) );
  INV_X1 U3518 ( .A(n3138), .ZN(n1066) );
  OAI22_X1 U3519 ( .A1(n3158), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[13][1] ), .B2(n3157), .ZN(n3139) );
  INV_X1 U3520 ( .A(n3139), .ZN(n1065) );
  OAI22_X1 U3521 ( .A1(n3158), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[13][2] ), .B2(n3157), .ZN(n3140) );
  INV_X1 U3522 ( .A(n3140), .ZN(n1064) );
  OAI22_X1 U3523 ( .A1(n3158), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[13][3] ), .B2(n3157), .ZN(n3141) );
  INV_X1 U3524 ( .A(n3141), .ZN(n1063) );
  OAI22_X1 U3525 ( .A1(n3158), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[13][4] ), .B2(n3157), .ZN(n3142) );
  INV_X1 U3526 ( .A(n3142), .ZN(n1062) );
  OAI22_X1 U3527 ( .A1(n3158), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[13][5] ), .B2(n3157), .ZN(n3143) );
  INV_X1 U3528 ( .A(n3143), .ZN(n1061) );
  OAI22_X1 U3529 ( .A1(n3158), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[13][6] ), .B2(n3157), .ZN(n3144) );
  INV_X1 U3530 ( .A(n3144), .ZN(n1060) );
  OAI22_X1 U3531 ( .A1(n3158), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[13][7] ), .B2(n3157), .ZN(n3145) );
  INV_X1 U3532 ( .A(n3145), .ZN(n1059) );
  OAI22_X1 U3533 ( .A1(n3158), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[13][8] ), .B2(n3157), .ZN(n3146) );
  INV_X1 U3534 ( .A(n3146), .ZN(n1058) );
  OAI22_X1 U3535 ( .A1(n3158), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[13][9] ), .B2(n3157), .ZN(n3147) );
  INV_X1 U3536 ( .A(n3147), .ZN(n1057) );
  OAI22_X1 U3537 ( .A1(n3158), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[13][10] ), .B2(n3157), .ZN(n3148) );
  INV_X1 U3538 ( .A(n3148), .ZN(n1056) );
  OAI22_X1 U3539 ( .A1(n3158), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[13][11] ), .B2(n3157), .ZN(n3149) );
  INV_X1 U3540 ( .A(n3149), .ZN(n1055) );
  OAI22_X1 U3541 ( .A1(n3158), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[13][12] ), .B2(n3157), .ZN(n3150) );
  INV_X1 U3542 ( .A(n3150), .ZN(n1054) );
  OAI22_X1 U3543 ( .A1(n3158), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[13][13] ), .B2(n3157), .ZN(n3151) );
  INV_X1 U3544 ( .A(n3151), .ZN(n1053) );
  OAI22_X1 U3545 ( .A1(n3158), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[13][14] ), .B2(n3157), .ZN(n3152) );
  INV_X1 U3546 ( .A(n3152), .ZN(n1052) );
  OAI22_X1 U3547 ( .A1(n3158), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[13][15] ), .B2(n3157), .ZN(n3153) );
  INV_X1 U3548 ( .A(n3153), .ZN(n1051) );
  OAI22_X1 U3549 ( .A1(n3158), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[13][16] ), .B2(n3157), .ZN(n3154) );
  INV_X1 U3550 ( .A(n3154), .ZN(n1050) );
  OAI22_X1 U3551 ( .A1(n3158), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[13][17] ), .B2(n3157), .ZN(n3155) );
  INV_X1 U3552 ( .A(n3155), .ZN(n1049) );
  OAI22_X1 U3553 ( .A1(n3158), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[13][18] ), .B2(n3157), .ZN(n3156) );
  INV_X1 U3554 ( .A(n3156), .ZN(n1048) );
  OAI22_X1 U3555 ( .A1(n3158), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[13][19] ), .B2(n3157), .ZN(n3159) );
  INV_X1 U3556 ( .A(n3159), .ZN(n1047) );
  OAI22_X1 U3557 ( .A1(n3181), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[14][0] ), .B2(n3180), .ZN(n3161) );
  INV_X1 U3558 ( .A(n3161), .ZN(n1046) );
  OAI22_X1 U3559 ( .A1(n3181), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[14][1] ), .B2(n3180), .ZN(n3162) );
  INV_X1 U3560 ( .A(n3162), .ZN(n1045) );
  OAI22_X1 U3561 ( .A1(n3181), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[14][2] ), .B2(n3180), .ZN(n3163) );
  INV_X1 U3562 ( .A(n3163), .ZN(n1044) );
  OAI22_X1 U3563 ( .A1(n3181), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[14][3] ), .B2(n3180), .ZN(n3164) );
  INV_X1 U3564 ( .A(n3164), .ZN(n1043) );
  OAI22_X1 U3565 ( .A1(n3181), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[14][4] ), .B2(n3180), .ZN(n3165) );
  INV_X1 U3566 ( .A(n3165), .ZN(n1042) );
  OAI22_X1 U3567 ( .A1(n3181), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[14][5] ), .B2(n3180), .ZN(n3166) );
  INV_X1 U3568 ( .A(n3166), .ZN(n1041) );
  OAI22_X1 U3569 ( .A1(n3181), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[14][6] ), .B2(n3180), .ZN(n3167) );
  INV_X1 U3570 ( .A(n3167), .ZN(n1040) );
  OAI22_X1 U3571 ( .A1(n3181), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[14][7] ), .B2(n3180), .ZN(n3168) );
  INV_X1 U3572 ( .A(n3168), .ZN(n1039) );
  OAI22_X1 U3573 ( .A1(n3181), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[14][8] ), .B2(n3180), .ZN(n3169) );
  INV_X1 U3574 ( .A(n3169), .ZN(n1038) );
  OAI22_X1 U3575 ( .A1(n3181), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[14][9] ), .B2(n3180), .ZN(n3170) );
  INV_X1 U3576 ( .A(n3170), .ZN(n1037) );
  OAI22_X1 U3577 ( .A1(n3181), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[14][10] ), .B2(n3180), .ZN(n3171) );
  INV_X1 U3578 ( .A(n3171), .ZN(n1036) );
  OAI22_X1 U3579 ( .A1(n3181), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[14][11] ), .B2(n3180), .ZN(n3172) );
  INV_X1 U3580 ( .A(n3172), .ZN(n1035) );
  OAI22_X1 U3581 ( .A1(n3181), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[14][12] ), .B2(n3180), .ZN(n3173) );
  INV_X1 U3582 ( .A(n3173), .ZN(n1034) );
  OAI22_X1 U3583 ( .A1(n3181), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[14][13] ), .B2(n3180), .ZN(n3174) );
  INV_X1 U3584 ( .A(n3174), .ZN(n1033) );
  OAI22_X1 U3585 ( .A1(n3181), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[14][14] ), .B2(n3180), .ZN(n3175) );
  INV_X1 U3586 ( .A(n3175), .ZN(n1032) );
  OAI22_X1 U3587 ( .A1(n3181), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[14][15] ), .B2(n3180), .ZN(n3176) );
  INV_X1 U3588 ( .A(n3176), .ZN(n1031) );
  OAI22_X1 U3589 ( .A1(n3181), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[14][16] ), .B2(n3180), .ZN(n3177) );
  INV_X1 U3590 ( .A(n3177), .ZN(n1030) );
  OAI22_X1 U3591 ( .A1(n3181), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[14][17] ), .B2(n3180), .ZN(n3178) );
  INV_X1 U3592 ( .A(n3178), .ZN(n1029) );
  OAI22_X1 U3593 ( .A1(n3181), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[14][18] ), .B2(n3180), .ZN(n3179) );
  INV_X1 U3594 ( .A(n3179), .ZN(n1028) );
  OAI22_X1 U3595 ( .A1(n3181), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[14][19] ), .B2(n3180), .ZN(n3182) );
  INV_X1 U3596 ( .A(n3182), .ZN(n1027) );
  OAI22_X1 U3597 ( .A1(n3205), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[15][0] ), .B2(n3204), .ZN(n3185) );
  INV_X1 U3598 ( .A(n3185), .ZN(n1026) );
  OAI22_X1 U3599 ( .A1(n3205), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[15][1] ), .B2(n3204), .ZN(n3186) );
  INV_X1 U3600 ( .A(n3186), .ZN(n1025) );
  OAI22_X1 U3601 ( .A1(n3205), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[15][2] ), .B2(n3204), .ZN(n3187) );
  INV_X1 U3602 ( .A(n3187), .ZN(n1024) );
  OAI22_X1 U3603 ( .A1(n3205), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[15][3] ), .B2(n3204), .ZN(n3188) );
  INV_X1 U3604 ( .A(n3188), .ZN(n1023) );
  OAI22_X1 U3605 ( .A1(n3205), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[15][4] ), .B2(n3204), .ZN(n3189) );
  INV_X1 U3606 ( .A(n3189), .ZN(n1022) );
  OAI22_X1 U3607 ( .A1(n3205), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[15][5] ), .B2(n3204), .ZN(n3190) );
  INV_X1 U3608 ( .A(n3190), .ZN(n1021) );
  OAI22_X1 U3609 ( .A1(n3205), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[15][6] ), .B2(n3204), .ZN(n3191) );
  INV_X1 U3610 ( .A(n3191), .ZN(n1020) );
  OAI22_X1 U3611 ( .A1(n3205), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[15][7] ), .B2(n3204), .ZN(n3192) );
  INV_X1 U3612 ( .A(n3192), .ZN(n1019) );
  OAI22_X1 U3613 ( .A1(n3205), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[15][8] ), .B2(n3204), .ZN(n3193) );
  INV_X1 U3614 ( .A(n3193), .ZN(n1018) );
  OAI22_X1 U3615 ( .A1(n3205), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[15][9] ), .B2(n3204), .ZN(n3194) );
  INV_X1 U3616 ( .A(n3194), .ZN(n1017) );
  OAI22_X1 U3617 ( .A1(n3205), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[15][10] ), .B2(n3204), .ZN(n3195) );
  INV_X1 U3618 ( .A(n3195), .ZN(n1016) );
  OAI22_X1 U3619 ( .A1(n3205), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[15][11] ), .B2(n3204), .ZN(n3196) );
  INV_X1 U3620 ( .A(n3196), .ZN(n1015) );
  OAI22_X1 U3621 ( .A1(n3205), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[15][12] ), .B2(n3204), .ZN(n3197) );
  INV_X1 U3622 ( .A(n3197), .ZN(n1014) );
  OAI22_X1 U3623 ( .A1(n3205), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[15][13] ), .B2(n3204), .ZN(n3198) );
  INV_X1 U3624 ( .A(n3198), .ZN(n1013) );
  OAI22_X1 U3625 ( .A1(n3205), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[15][14] ), .B2(n3204), .ZN(n3199) );
  INV_X1 U3626 ( .A(n3199), .ZN(n1012) );
  OAI22_X1 U3627 ( .A1(n3205), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[15][15] ), .B2(n3204), .ZN(n3200) );
  INV_X1 U3628 ( .A(n3200), .ZN(n1011) );
  OAI22_X1 U3629 ( .A1(n3205), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[15][16] ), .B2(n3204), .ZN(n3201) );
  INV_X1 U3630 ( .A(n3201), .ZN(n1010) );
  OAI22_X1 U3631 ( .A1(n3205), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[15][17] ), .B2(n3204), .ZN(n3202) );
  INV_X1 U3632 ( .A(n3202), .ZN(n1009) );
  OAI22_X1 U3633 ( .A1(n3205), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[15][18] ), .B2(n3204), .ZN(n3203) );
  INV_X1 U3634 ( .A(n3203), .ZN(n1008) );
  OAI22_X1 U3635 ( .A1(n3205), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[15][19] ), .B2(n3204), .ZN(n3206) );
  INV_X1 U3636 ( .A(n3206), .ZN(n1007) );
  OAI22_X1 U3637 ( .A1(n3228), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[16][0] ), .B2(n3227), .ZN(n3208) );
  INV_X1 U3638 ( .A(n3208), .ZN(n1006) );
  OAI22_X1 U3639 ( .A1(n3228), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[16][1] ), .B2(n3227), .ZN(n3209) );
  INV_X1 U3640 ( .A(n3209), .ZN(n1005) );
  OAI22_X1 U3641 ( .A1(n3228), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[16][2] ), .B2(n3227), .ZN(n3210) );
  INV_X1 U3642 ( .A(n3210), .ZN(n1004) );
  OAI22_X1 U3643 ( .A1(n3228), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[16][3] ), .B2(n3227), .ZN(n3211) );
  INV_X1 U3644 ( .A(n3211), .ZN(n1003) );
  OAI22_X1 U3645 ( .A1(n3228), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[16][4] ), .B2(n3227), .ZN(n3212) );
  INV_X1 U3646 ( .A(n3212), .ZN(n1002) );
  OAI22_X1 U3647 ( .A1(n3228), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[16][5] ), .B2(n3227), .ZN(n3213) );
  INV_X1 U3648 ( .A(n3213), .ZN(n1001) );
  OAI22_X1 U3649 ( .A1(n3228), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[16][6] ), .B2(n3227), .ZN(n3214) );
  INV_X1 U3650 ( .A(n3214), .ZN(n1000) );
  OAI22_X1 U3651 ( .A1(n3228), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[16][7] ), .B2(n3227), .ZN(n3215) );
  INV_X1 U3652 ( .A(n3215), .ZN(n999) );
  OAI22_X1 U3653 ( .A1(n3228), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[16][8] ), .B2(n3227), .ZN(n3216) );
  INV_X1 U3654 ( .A(n3216), .ZN(n998) );
  OAI22_X1 U3655 ( .A1(n3228), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[16][9] ), .B2(n3227), .ZN(n3217) );
  INV_X1 U3656 ( .A(n3217), .ZN(n997) );
  OAI22_X1 U3657 ( .A1(n3228), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[16][10] ), .B2(n3227), .ZN(n3218) );
  INV_X1 U3658 ( .A(n3218), .ZN(n996) );
  OAI22_X1 U3659 ( .A1(n3228), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[16][11] ), .B2(n3227), .ZN(n3219) );
  INV_X1 U3660 ( .A(n3219), .ZN(n995) );
  OAI22_X1 U3661 ( .A1(n3228), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[16][12] ), .B2(n3227), .ZN(n3220) );
  INV_X1 U3662 ( .A(n3220), .ZN(n994) );
  OAI22_X1 U3663 ( .A1(n3228), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[16][13] ), .B2(n3227), .ZN(n3221) );
  INV_X1 U3664 ( .A(n3221), .ZN(n993) );
  OAI22_X1 U3665 ( .A1(n3228), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[16][14] ), .B2(n3227), .ZN(n3222) );
  INV_X1 U3666 ( .A(n3222), .ZN(n992) );
  OAI22_X1 U3667 ( .A1(n3228), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[16][15] ), .B2(n3227), .ZN(n3223) );
  INV_X1 U3668 ( .A(n3223), .ZN(n991) );
  OAI22_X1 U3669 ( .A1(n3228), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[16][16] ), .B2(n3227), .ZN(n3224) );
  INV_X1 U3670 ( .A(n3224), .ZN(n990) );
  OAI22_X1 U3671 ( .A1(n3228), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[16][17] ), .B2(n3227), .ZN(n3225) );
  INV_X1 U3672 ( .A(n3225), .ZN(n989) );
  OAI22_X1 U3673 ( .A1(n3228), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[16][18] ), .B2(n3227), .ZN(n3226) );
  INV_X1 U3674 ( .A(n3226), .ZN(n988) );
  OAI22_X1 U3675 ( .A1(n3228), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[16][19] ), .B2(n3227), .ZN(n3229) );
  INV_X1 U3676 ( .A(n3229), .ZN(n987) );
  OAI22_X1 U3677 ( .A1(n3251), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[17][0] ), .B2(n3250), .ZN(n3231) );
  INV_X1 U3678 ( .A(n3231), .ZN(n986) );
  OAI22_X1 U3679 ( .A1(n3251), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[17][1] ), .B2(n3250), .ZN(n3232) );
  INV_X1 U3680 ( .A(n3232), .ZN(n985) );
  OAI22_X1 U3681 ( .A1(n3251), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[17][2] ), .B2(n3250), .ZN(n3233) );
  INV_X1 U3682 ( .A(n3233), .ZN(n984) );
  OAI22_X1 U3683 ( .A1(n3251), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[17][3] ), .B2(n3250), .ZN(n3234) );
  INV_X1 U3684 ( .A(n3234), .ZN(n983) );
  OAI22_X1 U3685 ( .A1(n3251), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[17][4] ), .B2(n3250), .ZN(n3235) );
  INV_X1 U3686 ( .A(n3235), .ZN(n982) );
  OAI22_X1 U3687 ( .A1(n3251), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[17][5] ), .B2(n3250), .ZN(n3236) );
  INV_X1 U3688 ( .A(n3236), .ZN(n981) );
  OAI22_X1 U3689 ( .A1(n3251), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[17][6] ), .B2(n3250), .ZN(n3237) );
  INV_X1 U3690 ( .A(n3237), .ZN(n980) );
  OAI22_X1 U3691 ( .A1(n3251), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[17][7] ), .B2(n3250), .ZN(n3238) );
  INV_X1 U3692 ( .A(n3238), .ZN(n979) );
  OAI22_X1 U3693 ( .A1(n3251), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[17][8] ), .B2(n3250), .ZN(n3239) );
  INV_X1 U3694 ( .A(n3239), .ZN(n978) );
  OAI22_X1 U3695 ( .A1(n3251), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[17][9] ), .B2(n3250), .ZN(n3240) );
  INV_X1 U3696 ( .A(n3240), .ZN(n977) );
  OAI22_X1 U3697 ( .A1(n3251), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[17][10] ), .B2(n3250), .ZN(n3241) );
  INV_X1 U3698 ( .A(n3241), .ZN(n976) );
  OAI22_X1 U3699 ( .A1(n3251), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[17][11] ), .B2(n3250), .ZN(n3242) );
  INV_X1 U3700 ( .A(n3242), .ZN(n975) );
  OAI22_X1 U3701 ( .A1(n3251), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[17][12] ), .B2(n3250), .ZN(n3243) );
  INV_X1 U3702 ( .A(n3243), .ZN(n974) );
  OAI22_X1 U3703 ( .A1(n3251), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[17][13] ), .B2(n3250), .ZN(n3244) );
  INV_X1 U3704 ( .A(n3244), .ZN(n973) );
  OAI22_X1 U3705 ( .A1(n3251), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[17][14] ), .B2(n3250), .ZN(n3245) );
  INV_X1 U3706 ( .A(n3245), .ZN(n972) );
  OAI22_X1 U3707 ( .A1(n3251), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[17][15] ), .B2(n3250), .ZN(n3246) );
  INV_X1 U3708 ( .A(n3246), .ZN(n971) );
  OAI22_X1 U3709 ( .A1(n3251), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[17][16] ), .B2(n3250), .ZN(n3247) );
  INV_X1 U3710 ( .A(n3247), .ZN(n970) );
  OAI22_X1 U3711 ( .A1(n3251), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[17][17] ), .B2(n3250), .ZN(n3248) );
  INV_X1 U3712 ( .A(n3248), .ZN(n969) );
  OAI22_X1 U3713 ( .A1(n3251), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[17][18] ), .B2(n3250), .ZN(n3249) );
  INV_X1 U3714 ( .A(n3249), .ZN(n968) );
  OAI22_X1 U3715 ( .A1(n3251), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[17][19] ), .B2(n3250), .ZN(n3252) );
  INV_X1 U3716 ( .A(n3252), .ZN(n967) );
  OAI22_X1 U3717 ( .A1(n3275), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[18][0] ), .B2(n3274), .ZN(n3255) );
  INV_X1 U3718 ( .A(n3255), .ZN(n966) );
  OAI22_X1 U3719 ( .A1(n3275), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[18][1] ), .B2(n3274), .ZN(n3256) );
  INV_X1 U3720 ( .A(n3256), .ZN(n965) );
  OAI22_X1 U3721 ( .A1(n3275), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[18][2] ), .B2(n3274), .ZN(n3257) );
  INV_X1 U3722 ( .A(n3257), .ZN(n964) );
  OAI22_X1 U3723 ( .A1(n3275), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[18][3] ), .B2(n3274), .ZN(n3258) );
  INV_X1 U3724 ( .A(n3258), .ZN(n963) );
  OAI22_X1 U3725 ( .A1(n3275), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[18][4] ), .B2(n3274), .ZN(n3259) );
  INV_X1 U3726 ( .A(n3259), .ZN(n962) );
  OAI22_X1 U3727 ( .A1(n3275), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[18][5] ), .B2(n3274), .ZN(n3260) );
  INV_X1 U3728 ( .A(n3260), .ZN(n961) );
  OAI22_X1 U3729 ( .A1(n3275), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[18][6] ), .B2(n3274), .ZN(n3261) );
  INV_X1 U3730 ( .A(n3261), .ZN(n960) );
  OAI22_X1 U3731 ( .A1(n3275), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[18][7] ), .B2(n3274), .ZN(n3262) );
  INV_X1 U3732 ( .A(n3262), .ZN(n959) );
  OAI22_X1 U3733 ( .A1(n3275), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[18][8] ), .B2(n3274), .ZN(n3263) );
  INV_X1 U3734 ( .A(n3263), .ZN(n958) );
  OAI22_X1 U3735 ( .A1(n3275), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[18][9] ), .B2(n3274), .ZN(n3264) );
  INV_X1 U3736 ( .A(n3264), .ZN(n957) );
  OAI22_X1 U3737 ( .A1(n3275), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[18][10] ), .B2(n3274), .ZN(n3265) );
  INV_X1 U3738 ( .A(n3265), .ZN(n956) );
  OAI22_X1 U3739 ( .A1(n3275), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[18][11] ), .B2(n3274), .ZN(n3266) );
  INV_X1 U3740 ( .A(n3266), .ZN(n955) );
  OAI22_X1 U3741 ( .A1(n3275), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[18][12] ), .B2(n3274), .ZN(n3267) );
  INV_X1 U3742 ( .A(n3267), .ZN(n954) );
  OAI22_X1 U3743 ( .A1(n3275), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[18][13] ), .B2(n3274), .ZN(n3268) );
  INV_X1 U3744 ( .A(n3268), .ZN(n953) );
  OAI22_X1 U3745 ( .A1(n3275), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[18][14] ), .B2(n3274), .ZN(n3269) );
  INV_X1 U3746 ( .A(n3269), .ZN(n952) );
  OAI22_X1 U3747 ( .A1(n3275), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[18][15] ), .B2(n3274), .ZN(n3270) );
  INV_X1 U3748 ( .A(n3270), .ZN(n951) );
  OAI22_X1 U3749 ( .A1(n3275), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[18][16] ), .B2(n3274), .ZN(n3271) );
  INV_X1 U3750 ( .A(n3271), .ZN(n950) );
  OAI22_X1 U3751 ( .A1(n3275), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[18][17] ), .B2(n3274), .ZN(n3272) );
  INV_X1 U3752 ( .A(n3272), .ZN(n949) );
  OAI22_X1 U3753 ( .A1(n3275), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[18][18] ), .B2(n3274), .ZN(n3273) );
  INV_X1 U3754 ( .A(n3273), .ZN(n948) );
  OAI22_X1 U3755 ( .A1(n3275), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[18][19] ), .B2(n3274), .ZN(n3276) );
  INV_X1 U3756 ( .A(n3276), .ZN(n947) );
  OAI22_X1 U3757 ( .A1(n3297), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[19][0] ), .B2(n3296), .ZN(n3277) );
  INV_X1 U3758 ( .A(n3277), .ZN(n946) );
  OAI22_X1 U3759 ( .A1(n3297), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[19][1] ), .B2(n3296), .ZN(n3278) );
  INV_X1 U3760 ( .A(n3278), .ZN(n945) );
  OAI22_X1 U3761 ( .A1(n3297), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[19][2] ), .B2(n3296), .ZN(n3279) );
  INV_X1 U3762 ( .A(n3279), .ZN(n944) );
  OAI22_X1 U3763 ( .A1(n3297), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[19][3] ), .B2(n3296), .ZN(n3280) );
  INV_X1 U3764 ( .A(n3280), .ZN(n943) );
  OAI22_X1 U3765 ( .A1(n3297), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[19][4] ), .B2(n3296), .ZN(n3281) );
  INV_X1 U3766 ( .A(n3281), .ZN(n942) );
  OAI22_X1 U3767 ( .A1(n3297), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[19][5] ), .B2(n3296), .ZN(n3282) );
  INV_X1 U3768 ( .A(n3282), .ZN(n941) );
  OAI22_X1 U3769 ( .A1(n3297), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[19][6] ), .B2(n3296), .ZN(n3283) );
  INV_X1 U3770 ( .A(n3283), .ZN(n940) );
  OAI22_X1 U3771 ( .A1(n3297), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[19][7] ), .B2(n3296), .ZN(n3284) );
  INV_X1 U3772 ( .A(n3284), .ZN(n939) );
  OAI22_X1 U3773 ( .A1(n3297), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[19][8] ), .B2(n3296), .ZN(n3285) );
  INV_X1 U3774 ( .A(n3285), .ZN(n938) );
  OAI22_X1 U3775 ( .A1(n3297), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[19][9] ), .B2(n3296), .ZN(n3286) );
  INV_X1 U3776 ( .A(n3286), .ZN(n937) );
  OAI22_X1 U3777 ( .A1(n3297), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[19][10] ), .B2(n3296), .ZN(n3287) );
  INV_X1 U3778 ( .A(n3287), .ZN(n936) );
  OAI22_X1 U3779 ( .A1(n3297), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[19][11] ), .B2(n3296), .ZN(n3288) );
  INV_X1 U3780 ( .A(n3288), .ZN(n935) );
  OAI22_X1 U3781 ( .A1(n3297), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[19][12] ), .B2(n3296), .ZN(n3289) );
  INV_X1 U3782 ( .A(n3289), .ZN(n934) );
  OAI22_X1 U3783 ( .A1(n3297), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[19][13] ), .B2(n3296), .ZN(n3290) );
  INV_X1 U3784 ( .A(n3290), .ZN(n933) );
  OAI22_X1 U3785 ( .A1(n3297), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[19][14] ), .B2(n3296), .ZN(n3291) );
  INV_X1 U3786 ( .A(n3291), .ZN(n932) );
  OAI22_X1 U3787 ( .A1(n3297), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[19][15] ), .B2(n3296), .ZN(n3292) );
  INV_X1 U3788 ( .A(n3292), .ZN(n931) );
  OAI22_X1 U3789 ( .A1(n3297), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[19][16] ), .B2(n3296), .ZN(n3293) );
  INV_X1 U3790 ( .A(n3293), .ZN(n930) );
  OAI22_X1 U3791 ( .A1(n3297), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[19][17] ), .B2(n3296), .ZN(n3294) );
  INV_X1 U3792 ( .A(n3294), .ZN(n929) );
  OAI22_X1 U3793 ( .A1(n3297), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[19][18] ), .B2(n3296), .ZN(n3295) );
  INV_X1 U3794 ( .A(n3295), .ZN(n928) );
  OAI22_X1 U3795 ( .A1(n3297), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[19][19] ), .B2(n3296), .ZN(n3298) );
  INV_X1 U3796 ( .A(n3298), .ZN(n927) );
  OAI22_X1 U3797 ( .A1(n3331), .A2(n3300), .B1(n3299), .B2(fmem_addr[0]), .ZN(
        n3301) );
  INV_X1 U3798 ( .A(n3301), .ZN(n926) );
  OAI222_X1 U3799 ( .A1(n3306), .A2(n3305), .B1(n3339), .B2(n3304), .C1(n3303), 
        .C2(n3302), .ZN(n923) );
  OAI22_X1 U3800 ( .A1(n3344), .A2(n3308), .B1(n3307), .B2(n3336), .ZN(n911)
         );
endmodule

