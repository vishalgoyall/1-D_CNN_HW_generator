
module conv_43_16_32_1 ( clk, reset, s_data_in_x, s_valid_x, s_ready_x, 
        m_data_out_y, m_valid_y, m_ready_y );
  input [31:0] s_data_in_x;
  output [31:0] m_data_out_y;
  input clk, reset, s_valid_x, m_ready_y;
  output s_ready_x, m_valid_y;
  wire   conv_done, conv_pre_start, N23, \fmem_inst/N78 , \fmem_inst/N77 ,
         \fmem_inst/N76 , \fmem_inst/N75 , \fmem_inst/N74 , \fmem_inst/N73 ,
         \fmem_inst/N72 , \fmem_inst/N71 , \fmem_inst/N70 , \fmem_inst/N69 ,
         \fmem_inst/N68 , \fmem_inst/N67 , \fmem_inst/N66 , \fmem_inst/N65 ,
         \fmem_inst/N64 , \fmem_inst/N63 , \fmem_inst/N62 ,
         \ctrl_conv_output_inst/N80 , \ctrl_conv_output_inst/N77 ,
         \ctrl_conv_output_inst/m_pre_valid_y ,
         \ctrl_conv_output_inst/conv_start_accum ,
         \ctrl_conv_output_inst/m_pre_pre_valid_y , n102, n103, n104, n105,
         n106, n107, n108, n109, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, \mac_unit_inst/n144 , \mac_unit_inst/n143 ,
         \mac_unit_inst/n142 , \mac_unit_inst/n141 , \mac_unit_inst/n140 ,
         \mac_unit_inst/n139 , \mac_unit_inst/n138 , \mac_unit_inst/n137 ,
         \mac_unit_inst/n136 , \mac_unit_inst/n135 , \mac_unit_inst/n134 ,
         \mac_unit_inst/n133 , \mac_unit_inst/n132 , \mac_unit_inst/n131 ,
         \mac_unit_inst/n130 , \mac_unit_inst/n129 , \mac_unit_inst/n128 ,
         \mac_unit_inst/n127 , \mac_unit_inst/n126 , \mac_unit_inst/n125 ,
         \mac_unit_inst/n124 , \mac_unit_inst/n123 , \mac_unit_inst/n122 ,
         \mac_unit_inst/n121 , \mac_unit_inst/n120 , \mac_unit_inst/n119 ,
         \mac_unit_inst/n118 , \mac_unit_inst/n117 , \mac_unit_inst/n116 ,
         \mac_unit_inst/n115 , \mac_unit_inst/n114 , \mac_unit_inst/n113 ,
         \mac_unit_inst/n112 , \mac_unit_inst/n111 , \mac_unit_inst/n110 ,
         \mac_unit_inst/n109 , \mac_unit_inst/n108 , \mac_unit_inst/n107 ,
         \mac_unit_inst/n106 , \mac_unit_inst/n105 , \mac_unit_inst/n104 ,
         \mac_unit_inst/n103 , \mac_unit_inst/n102 , \mac_unit_inst/n101 ,
         \mac_unit_inst/n100 , \mac_unit_inst/n99 , \mac_unit_inst/n98 ,
         \mac_unit_inst/n97 , \mac_unit_inst/n96 , \mac_unit_inst/n95 ,
         \mac_unit_inst/n94 , \mac_unit_inst/n93 , \mac_unit_inst/n92 ,
         \mac_unit_inst/n91 , \mac_unit_inst/n90 , \mac_unit_inst/n89 ,
         \mac_unit_inst/n88 , \mac_unit_inst/n87 , \mac_unit_inst/n86 ,
         \mac_unit_inst/n85 , \mac_unit_inst/n84 , \mac_unit_inst/n83 ,
         \mac_unit_inst/n82 , \mac_unit_inst/n81 , \xmem_inst/n3817 ,
         \xmem_inst/n3816 , \xmem_inst/n3815 , \xmem_inst/n3814 ,
         \xmem_inst/n3813 , \xmem_inst/n3812 , \xmem_inst/n3811 ,
         \xmem_inst/n3810 , \xmem_inst/n3809 , \xmem_inst/n3808 ,
         \xmem_inst/n3807 , \xmem_inst/n3806 , \xmem_inst/n3805 ,
         \xmem_inst/n3804 , \xmem_inst/n3803 , \xmem_inst/n3802 ,
         \xmem_inst/n3801 , \xmem_inst/n3800 , \xmem_inst/n3799 ,
         \xmem_inst/n3798 , \xmem_inst/n3797 , \xmem_inst/n3796 ,
         \xmem_inst/n3795 , \xmem_inst/n3794 , \xmem_inst/n3793 ,
         \xmem_inst/n3792 , \xmem_inst/n3791 , \xmem_inst/n3790 ,
         \xmem_inst/n3789 , \xmem_inst/n3788 , \xmem_inst/n3787 ,
         \xmem_inst/n3786 , \xmem_inst/n3785 , \xmem_inst/n3784 ,
         \xmem_inst/n3783 , \xmem_inst/n3782 , \xmem_inst/n3781 ,
         \xmem_inst/n3780 , \xmem_inst/n3779 , \xmem_inst/n3778 ,
         \xmem_inst/n3777 , \xmem_inst/n3776 , \xmem_inst/n3775 ,
         \xmem_inst/n3774 , \xmem_inst/n3773 , \xmem_inst/n3772 ,
         \xmem_inst/n3771 , \xmem_inst/n3770 , \xmem_inst/n3769 ,
         \xmem_inst/n3768 , \xmem_inst/n3767 , \xmem_inst/n3766 ,
         \xmem_inst/n3765 , \xmem_inst/n3764 , \xmem_inst/n3763 ,
         \xmem_inst/n3762 , \xmem_inst/n3761 , \xmem_inst/n3760 ,
         \xmem_inst/n3759 , \xmem_inst/n3758 , \xmem_inst/n3757 ,
         \xmem_inst/n3756 , \xmem_inst/n3755 , \xmem_inst/n3754 ,
         \xmem_inst/n3753 , \xmem_inst/n3752 , \xmem_inst/n3751 ,
         \xmem_inst/n3750 , \xmem_inst/n3749 , \xmem_inst/n3748 ,
         \xmem_inst/n3747 , \xmem_inst/n3746 , \xmem_inst/n3745 ,
         \xmem_inst/n3744 , \xmem_inst/n3743 , \xmem_inst/n3742 ,
         \xmem_inst/n3741 , \xmem_inst/n3740 , \xmem_inst/n3739 ,
         \xmem_inst/n3738 , \xmem_inst/n3737 , \xmem_inst/n3736 ,
         \xmem_inst/n3735 , \xmem_inst/n3734 , \xmem_inst/n3733 ,
         \xmem_inst/n3732 , \xmem_inst/n3731 , \xmem_inst/n3730 ,
         \xmem_inst/n3729 , \xmem_inst/n3728 , \xmem_inst/n3727 ,
         \xmem_inst/n3726 , \xmem_inst/n3725 , \xmem_inst/n3724 ,
         \xmem_inst/n3723 , \xmem_inst/n3722 , \xmem_inst/n3694 ,
         \xmem_inst/n3574 , \xmem_inst/n3559 , \xmem_inst/n3557 ,
         \xmem_inst/n3555 , \xmem_inst/n3544 , \xmem_inst/n3541 ,
         \xmem_inst/n3539 , \xmem_inst/n3538 , \xmem_inst/n3537 ,
         \xmem_inst/n3536 , \xmem_inst/n3535 , \xmem_inst/n3527 ,
         \xmem_inst/n3525 , \xmem_inst/n3523 , \xmem_inst/n3516 ,
         \xmem_inst/n3515 , \xmem_inst/n3514 , \xmem_inst/n3512 ,
         \xmem_inst/n3511 , \xmem_inst/n3510 , \xmem_inst/n3509 ,
         \xmem_inst/n3508 , \xmem_inst/n3507 , \xmem_inst/n3506 ,
         \xmem_inst/n3505 , \xmem_inst/n3504 , \xmem_inst/n3503 ,
         \xmem_inst/n3502 , \xmem_inst/n3501 , \xmem_inst/n3500 ,
         \xmem_inst/n3499 , \xmem_inst/n3498 , \xmem_inst/n3495 ,
         \xmem_inst/n3494 , \xmem_inst/n3493 , \xmem_inst/n3492 ,
         \xmem_inst/n3491 , \xmem_inst/n3490 , \xmem_inst/n3489 ,
         \xmem_inst/n3488 , \xmem_inst/n3487 , \xmem_inst/n3486 ,
         \xmem_inst/n3484 , \xmem_inst/n3483 , \xmem_inst/n3482 ,
         \xmem_inst/n3480 , \xmem_inst/n3479 , \xmem_inst/n3478 ,
         \xmem_inst/n3477 , \xmem_inst/n3476 , \xmem_inst/n3475 ,
         \xmem_inst/n3474 , \xmem_inst/n3473 , \xmem_inst/n3472 ,
         \xmem_inst/n3471 , \xmem_inst/n3470 , \xmem_inst/n3469 ,
         \xmem_inst/n3468 , \xmem_inst/n3467 , \xmem_inst/n3466 ,
         \xmem_inst/n2686 , \xmem_inst/N279 , \xmem_inst/N278 ,
         \xmem_inst/N277 , \xmem_inst/N276 , \xmem_inst/N275 ,
         \xmem_inst/N274 , \xmem_inst/N273 , \xmem_inst/N272 ,
         \xmem_inst/N271 , \xmem_inst/N270 , \xmem_inst/N269 ,
         \xmem_inst/N268 , \xmem_inst/N267 , \xmem_inst/N266 ,
         \xmem_inst/N265 , \xmem_inst/N264 , \xmem_inst/N263 ,
         \xmem_inst/N262 , \xmem_inst/N261 , \xmem_inst/N260 ,
         \xmem_inst/N259 , \xmem_inst/N258 , \xmem_inst/N257 ,
         \xmem_inst/N256 , \xmem_inst/N255 , \xmem_inst/N254 ,
         \xmem_inst/N253 , \xmem_inst/N252 , \xmem_inst/N251 ,
         \xmem_inst/N250 , \xmem_inst/N249 , \xmem_inst/N248 ,
         \xmem_inst/mem[42][31] , \xmem_inst/mem[42][30] ,
         \xmem_inst/mem[42][29] , \xmem_inst/mem[42][28] ,
         \xmem_inst/mem[42][27] , \xmem_inst/mem[42][26] ,
         \xmem_inst/mem[42][25] , \xmem_inst/mem[42][24] ,
         \xmem_inst/mem[42][23] , \xmem_inst/mem[42][22] ,
         \xmem_inst/mem[42][21] , \xmem_inst/mem[42][20] ,
         \xmem_inst/mem[42][19] , \xmem_inst/mem[42][18] ,
         \xmem_inst/mem[42][17] , \xmem_inst/mem[42][16] ,
         \xmem_inst/mem[42][15] , \xmem_inst/mem[42][14] ,
         \xmem_inst/mem[42][13] , \xmem_inst/mem[42][12] ,
         \xmem_inst/mem[42][11] , \xmem_inst/mem[42][10] ,
         \xmem_inst/mem[42][9] , \xmem_inst/mem[42][8] ,
         \xmem_inst/mem[42][7] , \xmem_inst/mem[42][6] ,
         \xmem_inst/mem[42][5] , \xmem_inst/mem[42][4] ,
         \xmem_inst/mem[42][3] , \xmem_inst/mem[42][2] ,
         \xmem_inst/mem[42][1] , \xmem_inst/mem[42][0] ,
         \xmem_inst/mem[41][31] , \xmem_inst/mem[41][30] ,
         \xmem_inst/mem[41][29] , \xmem_inst/mem[41][28] ,
         \xmem_inst/mem[41][27] , \xmem_inst/mem[41][26] ,
         \xmem_inst/mem[41][25] , \xmem_inst/mem[41][24] ,
         \xmem_inst/mem[41][23] , \xmem_inst/mem[41][22] ,
         \xmem_inst/mem[41][21] , \xmem_inst/mem[41][20] ,
         \xmem_inst/mem[41][19] , \xmem_inst/mem[41][18] ,
         \xmem_inst/mem[41][17] , \xmem_inst/mem[41][16] ,
         \xmem_inst/mem[41][15] , \xmem_inst/mem[41][14] ,
         \xmem_inst/mem[41][13] , \xmem_inst/mem[41][12] ,
         \xmem_inst/mem[41][11] , \xmem_inst/mem[41][10] ,
         \xmem_inst/mem[41][9] , \xmem_inst/mem[41][8] ,
         \xmem_inst/mem[41][7] , \xmem_inst/mem[41][6] ,
         \xmem_inst/mem[41][5] , \xmem_inst/mem[41][4] ,
         \xmem_inst/mem[41][3] , \xmem_inst/mem[41][2] ,
         \xmem_inst/mem[41][1] , \xmem_inst/mem[41][0] ,
         \xmem_inst/mem[40][31] , \xmem_inst/mem[40][30] ,
         \xmem_inst/mem[40][29] , \xmem_inst/mem[40][28] ,
         \xmem_inst/mem[40][27] , \xmem_inst/mem[40][26] ,
         \xmem_inst/mem[40][25] , \xmem_inst/mem[40][24] ,
         \xmem_inst/mem[40][23] , \xmem_inst/mem[40][22] ,
         \xmem_inst/mem[40][21] , \xmem_inst/mem[40][20] ,
         \xmem_inst/mem[40][19] , \xmem_inst/mem[40][18] ,
         \xmem_inst/mem[40][17] , \xmem_inst/mem[40][16] ,
         \xmem_inst/mem[40][15] , \xmem_inst/mem[40][14] ,
         \xmem_inst/mem[40][13] , \xmem_inst/mem[40][12] ,
         \xmem_inst/mem[40][11] , \xmem_inst/mem[40][10] ,
         \xmem_inst/mem[40][9] , \xmem_inst/mem[40][8] ,
         \xmem_inst/mem[40][7] , \xmem_inst/mem[40][6] ,
         \xmem_inst/mem[40][5] , \xmem_inst/mem[40][4] ,
         \xmem_inst/mem[40][3] , \xmem_inst/mem[40][2] ,
         \xmem_inst/mem[40][1] , \xmem_inst/mem[40][0] ,
         \xmem_inst/mem[39][31] , \xmem_inst/mem[39][30] ,
         \xmem_inst/mem[39][29] , \xmem_inst/mem[39][28] ,
         \xmem_inst/mem[39][27] , \xmem_inst/mem[39][26] ,
         \xmem_inst/mem[39][25] , \xmem_inst/mem[39][24] ,
         \xmem_inst/mem[39][23] , \xmem_inst/mem[39][22] ,
         \xmem_inst/mem[39][21] , \xmem_inst/mem[39][20] ,
         \xmem_inst/mem[39][19] , \xmem_inst/mem[39][18] ,
         \xmem_inst/mem[39][17] , \xmem_inst/mem[39][16] ,
         \xmem_inst/mem[39][15] , \xmem_inst/mem[39][14] ,
         \xmem_inst/mem[39][13] , \xmem_inst/mem[39][12] ,
         \xmem_inst/mem[39][11] , \xmem_inst/mem[39][10] ,
         \xmem_inst/mem[39][9] , \xmem_inst/mem[39][8] ,
         \xmem_inst/mem[39][7] , \xmem_inst/mem[39][6] ,
         \xmem_inst/mem[39][5] , \xmem_inst/mem[39][4] ,
         \xmem_inst/mem[39][3] , \xmem_inst/mem[39][2] ,
         \xmem_inst/mem[39][1] , \xmem_inst/mem[39][0] ,
         \xmem_inst/mem[38][31] , \xmem_inst/mem[38][30] ,
         \xmem_inst/mem[38][29] , \xmem_inst/mem[38][28] ,
         \xmem_inst/mem[38][27] , \xmem_inst/mem[38][26] ,
         \xmem_inst/mem[38][25] , \xmem_inst/mem[38][24] ,
         \xmem_inst/mem[38][23] , \xmem_inst/mem[38][22] ,
         \xmem_inst/mem[38][21] , \xmem_inst/mem[38][20] ,
         \xmem_inst/mem[38][19] , \xmem_inst/mem[38][18] ,
         \xmem_inst/mem[38][17] , \xmem_inst/mem[38][16] ,
         \xmem_inst/mem[38][15] , \xmem_inst/mem[38][14] ,
         \xmem_inst/mem[38][13] , \xmem_inst/mem[38][12] ,
         \xmem_inst/mem[38][11] , \xmem_inst/mem[38][10] ,
         \xmem_inst/mem[38][9] , \xmem_inst/mem[38][8] ,
         \xmem_inst/mem[38][7] , \xmem_inst/mem[38][6] ,
         \xmem_inst/mem[38][5] , \xmem_inst/mem[38][4] ,
         \xmem_inst/mem[38][3] , \xmem_inst/mem[38][2] ,
         \xmem_inst/mem[38][1] , \xmem_inst/mem[38][0] ,
         \xmem_inst/mem[37][31] , \xmem_inst/mem[37][30] ,
         \xmem_inst/mem[37][29] , \xmem_inst/mem[37][28] ,
         \xmem_inst/mem[37][27] , \xmem_inst/mem[37][26] ,
         \xmem_inst/mem[37][25] , \xmem_inst/mem[37][24] ,
         \xmem_inst/mem[37][23] , \xmem_inst/mem[37][22] ,
         \xmem_inst/mem[37][21] , \xmem_inst/mem[37][20] ,
         \xmem_inst/mem[37][19] , \xmem_inst/mem[37][18] ,
         \xmem_inst/mem[37][17] , \xmem_inst/mem[37][16] ,
         \xmem_inst/mem[37][15] , \xmem_inst/mem[37][14] ,
         \xmem_inst/mem[37][13] , \xmem_inst/mem[37][12] ,
         \xmem_inst/mem[37][11] , \xmem_inst/mem[37][10] ,
         \xmem_inst/mem[37][9] , \xmem_inst/mem[37][8] ,
         \xmem_inst/mem[37][7] , \xmem_inst/mem[37][6] ,
         \xmem_inst/mem[37][5] , \xmem_inst/mem[37][4] ,
         \xmem_inst/mem[37][3] , \xmem_inst/mem[37][2] ,
         \xmem_inst/mem[37][1] , \xmem_inst/mem[37][0] ,
         \xmem_inst/mem[36][31] , \xmem_inst/mem[36][30] ,
         \xmem_inst/mem[36][29] , \xmem_inst/mem[36][28] ,
         \xmem_inst/mem[36][27] , \xmem_inst/mem[36][26] ,
         \xmem_inst/mem[36][25] , \xmem_inst/mem[36][24] ,
         \xmem_inst/mem[36][23] , \xmem_inst/mem[36][22] ,
         \xmem_inst/mem[36][21] , \xmem_inst/mem[36][20] ,
         \xmem_inst/mem[36][19] , \xmem_inst/mem[36][18] ,
         \xmem_inst/mem[36][17] , \xmem_inst/mem[36][16] ,
         \xmem_inst/mem[36][15] , \xmem_inst/mem[36][14] ,
         \xmem_inst/mem[36][13] , \xmem_inst/mem[36][12] ,
         \xmem_inst/mem[36][11] , \xmem_inst/mem[36][10] ,
         \xmem_inst/mem[36][9] , \xmem_inst/mem[36][8] ,
         \xmem_inst/mem[36][7] , \xmem_inst/mem[36][6] ,
         \xmem_inst/mem[36][5] , \xmem_inst/mem[36][4] ,
         \xmem_inst/mem[36][3] , \xmem_inst/mem[36][2] ,
         \xmem_inst/mem[36][1] , \xmem_inst/mem[36][0] ,
         \xmem_inst/mem[35][31] , \xmem_inst/mem[35][30] ,
         \xmem_inst/mem[35][29] , \xmem_inst/mem[35][28] ,
         \xmem_inst/mem[35][27] , \xmem_inst/mem[35][26] ,
         \xmem_inst/mem[35][25] , \xmem_inst/mem[35][24] ,
         \xmem_inst/mem[35][23] , \xmem_inst/mem[35][22] ,
         \xmem_inst/mem[35][21] , \xmem_inst/mem[35][20] ,
         \xmem_inst/mem[35][19] , \xmem_inst/mem[35][18] ,
         \xmem_inst/mem[35][17] , \xmem_inst/mem[35][16] ,
         \xmem_inst/mem[35][15] , \xmem_inst/mem[35][14] ,
         \xmem_inst/mem[35][13] , \xmem_inst/mem[35][12] ,
         \xmem_inst/mem[35][11] , \xmem_inst/mem[35][10] ,
         \xmem_inst/mem[35][9] , \xmem_inst/mem[35][8] ,
         \xmem_inst/mem[35][7] , \xmem_inst/mem[35][6] ,
         \xmem_inst/mem[35][5] , \xmem_inst/mem[35][4] ,
         \xmem_inst/mem[35][3] , \xmem_inst/mem[35][2] ,
         \xmem_inst/mem[35][1] , \xmem_inst/mem[35][0] ,
         \xmem_inst/mem[34][31] , \xmem_inst/mem[34][30] ,
         \xmem_inst/mem[34][29] , \xmem_inst/mem[34][28] ,
         \xmem_inst/mem[34][27] , \xmem_inst/mem[34][26] ,
         \xmem_inst/mem[34][25] , \xmem_inst/mem[34][24] ,
         \xmem_inst/mem[34][23] , \xmem_inst/mem[34][22] ,
         \xmem_inst/mem[34][21] , \xmem_inst/mem[34][20] ,
         \xmem_inst/mem[34][19] , \xmem_inst/mem[34][18] ,
         \xmem_inst/mem[34][17] , \xmem_inst/mem[34][16] ,
         \xmem_inst/mem[34][15] , \xmem_inst/mem[34][14] ,
         \xmem_inst/mem[34][13] , \xmem_inst/mem[34][12] ,
         \xmem_inst/mem[34][11] , \xmem_inst/mem[34][10] ,
         \xmem_inst/mem[34][9] , \xmem_inst/mem[34][8] ,
         \xmem_inst/mem[34][7] , \xmem_inst/mem[34][6] ,
         \xmem_inst/mem[34][5] , \xmem_inst/mem[34][4] ,
         \xmem_inst/mem[34][3] , \xmem_inst/mem[34][2] ,
         \xmem_inst/mem[34][1] , \xmem_inst/mem[34][0] ,
         \xmem_inst/mem[33][31] , \xmem_inst/mem[33][30] ,
         \xmem_inst/mem[33][29] , \xmem_inst/mem[33][28] ,
         \xmem_inst/mem[33][27] , \xmem_inst/mem[33][26] ,
         \xmem_inst/mem[33][25] , \xmem_inst/mem[33][24] ,
         \xmem_inst/mem[33][23] , \xmem_inst/mem[33][22] ,
         \xmem_inst/mem[33][21] , \xmem_inst/mem[33][20] ,
         \xmem_inst/mem[33][19] , \xmem_inst/mem[33][18] ,
         \xmem_inst/mem[33][17] , \xmem_inst/mem[33][16] ,
         \xmem_inst/mem[33][15] , \xmem_inst/mem[33][14] ,
         \xmem_inst/mem[33][13] , \xmem_inst/mem[33][12] ,
         \xmem_inst/mem[33][11] , \xmem_inst/mem[33][10] ,
         \xmem_inst/mem[33][9] , \xmem_inst/mem[33][8] ,
         \xmem_inst/mem[33][7] , \xmem_inst/mem[33][6] ,
         \xmem_inst/mem[33][5] , \xmem_inst/mem[33][4] ,
         \xmem_inst/mem[33][3] , \xmem_inst/mem[33][2] ,
         \xmem_inst/mem[33][1] , \xmem_inst/mem[33][0] ,
         \xmem_inst/mem[32][31] , \xmem_inst/mem[32][30] ,
         \xmem_inst/mem[32][29] , \xmem_inst/mem[32][28] ,
         \xmem_inst/mem[32][27] , \xmem_inst/mem[32][26] ,
         \xmem_inst/mem[32][25] , \xmem_inst/mem[32][24] ,
         \xmem_inst/mem[32][23] , \xmem_inst/mem[32][22] ,
         \xmem_inst/mem[32][21] , \xmem_inst/mem[32][20] ,
         \xmem_inst/mem[32][19] , \xmem_inst/mem[32][18] ,
         \xmem_inst/mem[32][17] , \xmem_inst/mem[32][16] ,
         \xmem_inst/mem[32][15] , \xmem_inst/mem[32][14] ,
         \xmem_inst/mem[32][13] , \xmem_inst/mem[32][12] ,
         \xmem_inst/mem[32][11] , \xmem_inst/mem[32][10] ,
         \xmem_inst/mem[32][9] , \xmem_inst/mem[32][8] ,
         \xmem_inst/mem[32][7] , \xmem_inst/mem[32][6] ,
         \xmem_inst/mem[32][5] , \xmem_inst/mem[32][4] ,
         \xmem_inst/mem[32][3] , \xmem_inst/mem[32][2] ,
         \xmem_inst/mem[32][1] , \xmem_inst/mem[32][0] ,
         \xmem_inst/mem[31][31] , \xmem_inst/mem[31][30] ,
         \xmem_inst/mem[31][29] , \xmem_inst/mem[31][28] ,
         \xmem_inst/mem[31][27] , \xmem_inst/mem[31][26] ,
         \xmem_inst/mem[31][25] , \xmem_inst/mem[31][24] ,
         \xmem_inst/mem[31][23] , \xmem_inst/mem[31][22] ,
         \xmem_inst/mem[31][21] , \xmem_inst/mem[31][20] ,
         \xmem_inst/mem[31][19] , \xmem_inst/mem[31][18] ,
         \xmem_inst/mem[31][17] , \xmem_inst/mem[31][16] ,
         \xmem_inst/mem[31][15] , \xmem_inst/mem[31][14] ,
         \xmem_inst/mem[31][13] , \xmem_inst/mem[31][12] ,
         \xmem_inst/mem[31][11] , \xmem_inst/mem[31][10] ,
         \xmem_inst/mem[31][9] , \xmem_inst/mem[31][8] ,
         \xmem_inst/mem[31][7] , \xmem_inst/mem[31][6] ,
         \xmem_inst/mem[31][5] , \xmem_inst/mem[31][4] ,
         \xmem_inst/mem[31][3] , \xmem_inst/mem[31][2] ,
         \xmem_inst/mem[31][1] , \xmem_inst/mem[31][0] ,
         \xmem_inst/mem[30][31] , \xmem_inst/mem[30][30] ,
         \xmem_inst/mem[30][29] , \xmem_inst/mem[30][28] ,
         \xmem_inst/mem[30][27] , \xmem_inst/mem[30][26] ,
         \xmem_inst/mem[30][25] , \xmem_inst/mem[30][24] ,
         \xmem_inst/mem[30][23] , \xmem_inst/mem[30][22] ,
         \xmem_inst/mem[30][21] , \xmem_inst/mem[30][20] ,
         \xmem_inst/mem[30][19] , \xmem_inst/mem[30][18] ,
         \xmem_inst/mem[30][17] , \xmem_inst/mem[30][16] ,
         \xmem_inst/mem[30][15] , \xmem_inst/mem[30][14] ,
         \xmem_inst/mem[30][13] , \xmem_inst/mem[30][12] ,
         \xmem_inst/mem[30][11] , \xmem_inst/mem[30][10] ,
         \xmem_inst/mem[30][9] , \xmem_inst/mem[30][8] ,
         \xmem_inst/mem[30][7] , \xmem_inst/mem[30][6] ,
         \xmem_inst/mem[30][5] , \xmem_inst/mem[30][4] ,
         \xmem_inst/mem[30][3] , \xmem_inst/mem[30][2] ,
         \xmem_inst/mem[30][1] , \xmem_inst/mem[30][0] ,
         \xmem_inst/mem[29][31] , \xmem_inst/mem[29][30] ,
         \xmem_inst/mem[29][29] , \xmem_inst/mem[29][28] ,
         \xmem_inst/mem[29][27] , \xmem_inst/mem[29][26] ,
         \xmem_inst/mem[29][25] , \xmem_inst/mem[29][24] ,
         \xmem_inst/mem[29][23] , \xmem_inst/mem[29][22] ,
         \xmem_inst/mem[29][21] , \xmem_inst/mem[29][20] ,
         \xmem_inst/mem[29][19] , \xmem_inst/mem[29][18] ,
         \xmem_inst/mem[29][17] , \xmem_inst/mem[29][16] ,
         \xmem_inst/mem[29][15] , \xmem_inst/mem[29][14] ,
         \xmem_inst/mem[29][13] , \xmem_inst/mem[29][12] ,
         \xmem_inst/mem[29][11] , \xmem_inst/mem[29][10] ,
         \xmem_inst/mem[29][9] , \xmem_inst/mem[29][8] ,
         \xmem_inst/mem[29][7] , \xmem_inst/mem[29][6] ,
         \xmem_inst/mem[29][5] , \xmem_inst/mem[29][4] ,
         \xmem_inst/mem[29][3] , \xmem_inst/mem[29][2] ,
         \xmem_inst/mem[29][1] , \xmem_inst/mem[29][0] ,
         \xmem_inst/mem[28][31] , \xmem_inst/mem[28][30] ,
         \xmem_inst/mem[28][29] , \xmem_inst/mem[28][28] ,
         \xmem_inst/mem[28][27] , \xmem_inst/mem[28][26] ,
         \xmem_inst/mem[28][25] , \xmem_inst/mem[28][24] ,
         \xmem_inst/mem[28][23] , \xmem_inst/mem[28][22] ,
         \xmem_inst/mem[28][21] , \xmem_inst/mem[28][20] ,
         \xmem_inst/mem[28][19] , \xmem_inst/mem[28][18] ,
         \xmem_inst/mem[28][17] , \xmem_inst/mem[28][16] ,
         \xmem_inst/mem[28][15] , \xmem_inst/mem[28][14] ,
         \xmem_inst/mem[28][13] , \xmem_inst/mem[28][12] ,
         \xmem_inst/mem[28][11] , \xmem_inst/mem[28][10] ,
         \xmem_inst/mem[28][9] , \xmem_inst/mem[28][8] ,
         \xmem_inst/mem[28][7] , \xmem_inst/mem[28][6] ,
         \xmem_inst/mem[28][5] , \xmem_inst/mem[28][4] ,
         \xmem_inst/mem[28][3] , \xmem_inst/mem[28][2] ,
         \xmem_inst/mem[28][1] , \xmem_inst/mem[28][0] ,
         \xmem_inst/mem[27][31] , \xmem_inst/mem[27][30] ,
         \xmem_inst/mem[27][29] , \xmem_inst/mem[27][28] ,
         \xmem_inst/mem[27][27] , \xmem_inst/mem[27][26] ,
         \xmem_inst/mem[27][25] , \xmem_inst/mem[27][24] ,
         \xmem_inst/mem[27][23] , \xmem_inst/mem[27][22] ,
         \xmem_inst/mem[27][21] , \xmem_inst/mem[27][20] ,
         \xmem_inst/mem[27][19] , \xmem_inst/mem[27][18] ,
         \xmem_inst/mem[27][17] , \xmem_inst/mem[27][16] ,
         \xmem_inst/mem[27][15] , \xmem_inst/mem[27][14] ,
         \xmem_inst/mem[27][13] , \xmem_inst/mem[27][12] ,
         \xmem_inst/mem[27][11] , \xmem_inst/mem[27][10] ,
         \xmem_inst/mem[27][9] , \xmem_inst/mem[27][8] ,
         \xmem_inst/mem[27][7] , \xmem_inst/mem[27][6] ,
         \xmem_inst/mem[27][5] , \xmem_inst/mem[27][4] ,
         \xmem_inst/mem[27][3] , \xmem_inst/mem[27][2] ,
         \xmem_inst/mem[27][1] , \xmem_inst/mem[27][0] ,
         \xmem_inst/mem[26][31] , \xmem_inst/mem[26][30] ,
         \xmem_inst/mem[26][29] , \xmem_inst/mem[26][28] ,
         \xmem_inst/mem[26][27] , \xmem_inst/mem[26][26] ,
         \xmem_inst/mem[26][25] , \xmem_inst/mem[26][24] ,
         \xmem_inst/mem[26][23] , \xmem_inst/mem[26][22] ,
         \xmem_inst/mem[26][21] , \xmem_inst/mem[26][20] ,
         \xmem_inst/mem[26][19] , \xmem_inst/mem[26][18] ,
         \xmem_inst/mem[26][17] , \xmem_inst/mem[26][16] ,
         \xmem_inst/mem[26][15] , \xmem_inst/mem[26][14] ,
         \xmem_inst/mem[26][13] , \xmem_inst/mem[26][12] ,
         \xmem_inst/mem[26][11] , \xmem_inst/mem[26][10] ,
         \xmem_inst/mem[26][9] , \xmem_inst/mem[26][8] ,
         \xmem_inst/mem[26][7] , \xmem_inst/mem[26][6] ,
         \xmem_inst/mem[26][5] , \xmem_inst/mem[26][4] ,
         \xmem_inst/mem[26][3] , \xmem_inst/mem[26][2] ,
         \xmem_inst/mem[26][1] , \xmem_inst/mem[26][0] ,
         \xmem_inst/mem[25][31] , \xmem_inst/mem[25][30] ,
         \xmem_inst/mem[25][29] , \xmem_inst/mem[25][28] ,
         \xmem_inst/mem[25][27] , \xmem_inst/mem[25][26] ,
         \xmem_inst/mem[25][25] , \xmem_inst/mem[25][24] ,
         \xmem_inst/mem[25][23] , \xmem_inst/mem[25][22] ,
         \xmem_inst/mem[25][21] , \xmem_inst/mem[25][20] ,
         \xmem_inst/mem[25][19] , \xmem_inst/mem[25][18] ,
         \xmem_inst/mem[25][17] , \xmem_inst/mem[25][16] ,
         \xmem_inst/mem[25][15] , \xmem_inst/mem[25][14] ,
         \xmem_inst/mem[25][13] , \xmem_inst/mem[25][12] ,
         \xmem_inst/mem[25][11] , \xmem_inst/mem[25][10] ,
         \xmem_inst/mem[25][9] , \xmem_inst/mem[25][8] ,
         \xmem_inst/mem[25][7] , \xmem_inst/mem[25][6] ,
         \xmem_inst/mem[25][5] , \xmem_inst/mem[25][4] ,
         \xmem_inst/mem[25][3] , \xmem_inst/mem[25][2] ,
         \xmem_inst/mem[25][1] , \xmem_inst/mem[25][0] ,
         \xmem_inst/mem[24][31] , \xmem_inst/mem[24][30] ,
         \xmem_inst/mem[24][29] , \xmem_inst/mem[24][28] ,
         \xmem_inst/mem[24][27] , \xmem_inst/mem[24][26] ,
         \xmem_inst/mem[24][25] , \xmem_inst/mem[24][24] ,
         \xmem_inst/mem[24][23] , \xmem_inst/mem[24][22] ,
         \xmem_inst/mem[24][21] , \xmem_inst/mem[24][20] ,
         \xmem_inst/mem[24][19] , \xmem_inst/mem[24][18] ,
         \xmem_inst/mem[24][17] , \xmem_inst/mem[24][16] ,
         \xmem_inst/mem[24][15] , \xmem_inst/mem[24][14] ,
         \xmem_inst/mem[24][13] , \xmem_inst/mem[24][12] ,
         \xmem_inst/mem[24][11] , \xmem_inst/mem[24][10] ,
         \xmem_inst/mem[24][9] , \xmem_inst/mem[24][8] ,
         \xmem_inst/mem[24][7] , \xmem_inst/mem[24][6] ,
         \xmem_inst/mem[24][5] , \xmem_inst/mem[24][4] ,
         \xmem_inst/mem[24][3] , \xmem_inst/mem[24][2] ,
         \xmem_inst/mem[24][1] , \xmem_inst/mem[24][0] ,
         \xmem_inst/mem[23][31] , \xmem_inst/mem[23][30] ,
         \xmem_inst/mem[23][29] , \xmem_inst/mem[23][28] ,
         \xmem_inst/mem[23][27] , \xmem_inst/mem[23][26] ,
         \xmem_inst/mem[23][25] , \xmem_inst/mem[23][24] ,
         \xmem_inst/mem[23][23] , \xmem_inst/mem[23][22] ,
         \xmem_inst/mem[23][21] , \xmem_inst/mem[23][20] ,
         \xmem_inst/mem[23][19] , \xmem_inst/mem[23][18] ,
         \xmem_inst/mem[23][17] , \xmem_inst/mem[23][16] ,
         \xmem_inst/mem[23][15] , \xmem_inst/mem[23][14] ,
         \xmem_inst/mem[23][13] , \xmem_inst/mem[23][12] ,
         \xmem_inst/mem[23][11] , \xmem_inst/mem[23][10] ,
         \xmem_inst/mem[23][9] , \xmem_inst/mem[23][8] ,
         \xmem_inst/mem[23][7] , \xmem_inst/mem[23][6] ,
         \xmem_inst/mem[23][5] , \xmem_inst/mem[23][4] ,
         \xmem_inst/mem[23][3] , \xmem_inst/mem[23][2] ,
         \xmem_inst/mem[23][1] , \xmem_inst/mem[23][0] ,
         \xmem_inst/mem[22][31] , \xmem_inst/mem[22][30] ,
         \xmem_inst/mem[22][29] , \xmem_inst/mem[22][28] ,
         \xmem_inst/mem[22][27] , \xmem_inst/mem[22][26] ,
         \xmem_inst/mem[22][25] , \xmem_inst/mem[22][24] ,
         \xmem_inst/mem[22][23] , \xmem_inst/mem[22][22] ,
         \xmem_inst/mem[22][21] , \xmem_inst/mem[22][20] ,
         \xmem_inst/mem[22][19] , \xmem_inst/mem[22][18] ,
         \xmem_inst/mem[22][17] , \xmem_inst/mem[22][16] ,
         \xmem_inst/mem[22][15] , \xmem_inst/mem[22][14] ,
         \xmem_inst/mem[22][13] , \xmem_inst/mem[22][12] ,
         \xmem_inst/mem[22][11] , \xmem_inst/mem[22][10] ,
         \xmem_inst/mem[22][9] , \xmem_inst/mem[22][8] ,
         \xmem_inst/mem[22][7] , \xmem_inst/mem[22][6] ,
         \xmem_inst/mem[22][5] , \xmem_inst/mem[22][4] ,
         \xmem_inst/mem[22][3] , \xmem_inst/mem[22][2] ,
         \xmem_inst/mem[22][1] , \xmem_inst/mem[22][0] ,
         \xmem_inst/mem[21][31] , \xmem_inst/mem[21][30] ,
         \xmem_inst/mem[21][29] , \xmem_inst/mem[21][28] ,
         \xmem_inst/mem[21][27] , \xmem_inst/mem[21][26] ,
         \xmem_inst/mem[21][25] , \xmem_inst/mem[21][24] ,
         \xmem_inst/mem[21][23] , \xmem_inst/mem[21][22] ,
         \xmem_inst/mem[21][21] , \xmem_inst/mem[21][20] ,
         \xmem_inst/mem[21][19] , \xmem_inst/mem[21][18] ,
         \xmem_inst/mem[21][17] , \xmem_inst/mem[21][16] ,
         \xmem_inst/mem[21][15] , \xmem_inst/mem[21][14] ,
         \xmem_inst/mem[21][13] , \xmem_inst/mem[21][12] ,
         \xmem_inst/mem[21][11] , \xmem_inst/mem[21][10] ,
         \xmem_inst/mem[21][9] , \xmem_inst/mem[21][8] ,
         \xmem_inst/mem[21][7] , \xmem_inst/mem[21][6] ,
         \xmem_inst/mem[21][5] , \xmem_inst/mem[21][4] ,
         \xmem_inst/mem[21][3] , \xmem_inst/mem[21][2] ,
         \xmem_inst/mem[21][1] , \xmem_inst/mem[21][0] ,
         \xmem_inst/mem[20][31] , \xmem_inst/mem[20][30] ,
         \xmem_inst/mem[20][29] , \xmem_inst/mem[20][28] ,
         \xmem_inst/mem[20][27] , \xmem_inst/mem[20][26] ,
         \xmem_inst/mem[20][25] , \xmem_inst/mem[20][24] ,
         \xmem_inst/mem[20][23] , \xmem_inst/mem[20][22] ,
         \xmem_inst/mem[20][21] , \xmem_inst/mem[20][20] ,
         \xmem_inst/mem[20][19] , \xmem_inst/mem[20][18] ,
         \xmem_inst/mem[20][17] , \xmem_inst/mem[20][16] ,
         \xmem_inst/mem[20][15] , \xmem_inst/mem[20][14] ,
         \xmem_inst/mem[20][13] , \xmem_inst/mem[20][12] ,
         \xmem_inst/mem[20][11] , \xmem_inst/mem[20][10] ,
         \xmem_inst/mem[20][9] , \xmem_inst/mem[20][8] ,
         \xmem_inst/mem[20][7] , \xmem_inst/mem[20][6] ,
         \xmem_inst/mem[20][5] , \xmem_inst/mem[20][4] ,
         \xmem_inst/mem[20][3] , \xmem_inst/mem[20][2] ,
         \xmem_inst/mem[20][1] , \xmem_inst/mem[20][0] ,
         \xmem_inst/mem[19][31] , \xmem_inst/mem[19][30] ,
         \xmem_inst/mem[19][29] , \xmem_inst/mem[19][28] ,
         \xmem_inst/mem[19][27] , \xmem_inst/mem[19][26] ,
         \xmem_inst/mem[19][25] , \xmem_inst/mem[19][24] ,
         \xmem_inst/mem[19][23] , \xmem_inst/mem[19][22] ,
         \xmem_inst/mem[19][21] , \xmem_inst/mem[19][20] ,
         \xmem_inst/mem[19][19] , \xmem_inst/mem[19][18] ,
         \xmem_inst/mem[19][17] , \xmem_inst/mem[19][16] ,
         \xmem_inst/mem[19][15] , \xmem_inst/mem[19][14] ,
         \xmem_inst/mem[19][13] , \xmem_inst/mem[19][12] ,
         \xmem_inst/mem[19][11] , \xmem_inst/mem[19][10] ,
         \xmem_inst/mem[19][9] , \xmem_inst/mem[19][8] ,
         \xmem_inst/mem[19][7] , \xmem_inst/mem[19][6] ,
         \xmem_inst/mem[19][5] , \xmem_inst/mem[19][4] ,
         \xmem_inst/mem[19][3] , \xmem_inst/mem[19][2] ,
         \xmem_inst/mem[19][1] , \xmem_inst/mem[19][0] ,
         \xmem_inst/mem[18][31] , \xmem_inst/mem[18][30] ,
         \xmem_inst/mem[18][29] , \xmem_inst/mem[18][28] ,
         \xmem_inst/mem[18][27] , \xmem_inst/mem[18][26] ,
         \xmem_inst/mem[18][25] , \xmem_inst/mem[18][24] ,
         \xmem_inst/mem[18][23] , \xmem_inst/mem[18][22] ,
         \xmem_inst/mem[18][21] , \xmem_inst/mem[18][20] ,
         \xmem_inst/mem[18][19] , \xmem_inst/mem[18][18] ,
         \xmem_inst/mem[18][17] , \xmem_inst/mem[18][16] ,
         \xmem_inst/mem[18][15] , \xmem_inst/mem[18][14] ,
         \xmem_inst/mem[18][13] , \xmem_inst/mem[18][12] ,
         \xmem_inst/mem[18][11] , \xmem_inst/mem[18][10] ,
         \xmem_inst/mem[18][9] , \xmem_inst/mem[18][8] ,
         \xmem_inst/mem[18][7] , \xmem_inst/mem[18][6] ,
         \xmem_inst/mem[18][5] , \xmem_inst/mem[18][4] ,
         \xmem_inst/mem[18][3] , \xmem_inst/mem[18][2] ,
         \xmem_inst/mem[18][1] , \xmem_inst/mem[18][0] ,
         \xmem_inst/mem[17][31] , \xmem_inst/mem[17][30] ,
         \xmem_inst/mem[17][29] , \xmem_inst/mem[17][28] ,
         \xmem_inst/mem[17][27] , \xmem_inst/mem[17][26] ,
         \xmem_inst/mem[17][25] , \xmem_inst/mem[17][24] ,
         \xmem_inst/mem[17][23] , \xmem_inst/mem[17][22] ,
         \xmem_inst/mem[17][21] , \xmem_inst/mem[17][20] ,
         \xmem_inst/mem[17][19] , \xmem_inst/mem[17][18] ,
         \xmem_inst/mem[17][17] , \xmem_inst/mem[17][16] ,
         \xmem_inst/mem[17][15] , \xmem_inst/mem[17][14] ,
         \xmem_inst/mem[17][13] , \xmem_inst/mem[17][12] ,
         \xmem_inst/mem[17][11] , \xmem_inst/mem[17][10] ,
         \xmem_inst/mem[17][9] , \xmem_inst/mem[17][8] ,
         \xmem_inst/mem[17][7] , \xmem_inst/mem[17][6] ,
         \xmem_inst/mem[17][5] , \xmem_inst/mem[17][4] ,
         \xmem_inst/mem[17][3] , \xmem_inst/mem[17][2] ,
         \xmem_inst/mem[17][1] , \xmem_inst/mem[17][0] ,
         \xmem_inst/mem[16][31] , \xmem_inst/mem[16][30] ,
         \xmem_inst/mem[16][29] , \xmem_inst/mem[16][28] ,
         \xmem_inst/mem[16][27] , \xmem_inst/mem[16][26] ,
         \xmem_inst/mem[16][25] , \xmem_inst/mem[16][24] ,
         \xmem_inst/mem[16][23] , \xmem_inst/mem[16][22] ,
         \xmem_inst/mem[16][21] , \xmem_inst/mem[16][20] ,
         \xmem_inst/mem[16][19] , \xmem_inst/mem[16][18] ,
         \xmem_inst/mem[16][17] , \xmem_inst/mem[16][16] ,
         \xmem_inst/mem[16][15] , \xmem_inst/mem[16][14] ,
         \xmem_inst/mem[16][13] , \xmem_inst/mem[16][12] ,
         \xmem_inst/mem[16][11] , \xmem_inst/mem[16][10] ,
         \xmem_inst/mem[16][9] , \xmem_inst/mem[16][8] ,
         \xmem_inst/mem[16][7] , \xmem_inst/mem[16][6] ,
         \xmem_inst/mem[16][5] , \xmem_inst/mem[16][4] ,
         \xmem_inst/mem[16][3] , \xmem_inst/mem[16][2] ,
         \xmem_inst/mem[16][1] , \xmem_inst/mem[16][0] ,
         \xmem_inst/mem[15][31] , \xmem_inst/mem[15][30] ,
         \xmem_inst/mem[15][29] , \xmem_inst/mem[15][28] ,
         \xmem_inst/mem[15][27] , \xmem_inst/mem[15][26] ,
         \xmem_inst/mem[15][25] , \xmem_inst/mem[15][24] ,
         \xmem_inst/mem[15][23] , \xmem_inst/mem[15][22] ,
         \xmem_inst/mem[15][21] , \xmem_inst/mem[15][20] ,
         \xmem_inst/mem[15][19] , \xmem_inst/mem[15][18] ,
         \xmem_inst/mem[15][17] , \xmem_inst/mem[15][16] ,
         \xmem_inst/mem[15][15] , \xmem_inst/mem[15][14] ,
         \xmem_inst/mem[15][13] , \xmem_inst/mem[15][12] ,
         \xmem_inst/mem[15][11] , \xmem_inst/mem[15][10] ,
         \xmem_inst/mem[15][9] , \xmem_inst/mem[15][8] ,
         \xmem_inst/mem[15][7] , \xmem_inst/mem[15][6] ,
         \xmem_inst/mem[15][5] , \xmem_inst/mem[15][4] ,
         \xmem_inst/mem[15][3] , \xmem_inst/mem[15][2] ,
         \xmem_inst/mem[15][1] , \xmem_inst/mem[15][0] ,
         \xmem_inst/mem[14][31] , \xmem_inst/mem[14][30] ,
         \xmem_inst/mem[14][29] , \xmem_inst/mem[14][28] ,
         \xmem_inst/mem[14][27] , \xmem_inst/mem[14][26] ,
         \xmem_inst/mem[14][25] , \xmem_inst/mem[14][24] ,
         \xmem_inst/mem[14][23] , \xmem_inst/mem[14][22] ,
         \xmem_inst/mem[14][21] , \xmem_inst/mem[14][20] ,
         \xmem_inst/mem[14][19] , \xmem_inst/mem[14][18] ,
         \xmem_inst/mem[14][17] , \xmem_inst/mem[14][16] ,
         \xmem_inst/mem[14][15] , \xmem_inst/mem[14][14] ,
         \xmem_inst/mem[14][13] , \xmem_inst/mem[14][12] ,
         \xmem_inst/mem[14][11] , \xmem_inst/mem[14][10] ,
         \xmem_inst/mem[14][9] , \xmem_inst/mem[14][8] ,
         \xmem_inst/mem[14][7] , \xmem_inst/mem[14][6] ,
         \xmem_inst/mem[14][5] , \xmem_inst/mem[14][4] ,
         \xmem_inst/mem[14][3] , \xmem_inst/mem[14][2] ,
         \xmem_inst/mem[14][1] , \xmem_inst/mem[14][0] ,
         \xmem_inst/mem[13][31] , \xmem_inst/mem[13][30] ,
         \xmem_inst/mem[13][29] , \xmem_inst/mem[13][28] ,
         \xmem_inst/mem[13][27] , \xmem_inst/mem[13][26] ,
         \xmem_inst/mem[13][25] , \xmem_inst/mem[13][24] ,
         \xmem_inst/mem[13][23] , \xmem_inst/mem[13][22] ,
         \xmem_inst/mem[13][21] , \xmem_inst/mem[13][20] ,
         \xmem_inst/mem[13][19] , \xmem_inst/mem[13][18] ,
         \xmem_inst/mem[13][17] , \xmem_inst/mem[13][16] ,
         \xmem_inst/mem[13][15] , \xmem_inst/mem[13][14] ,
         \xmem_inst/mem[13][13] , \xmem_inst/mem[13][12] ,
         \xmem_inst/mem[13][11] , \xmem_inst/mem[13][10] ,
         \xmem_inst/mem[13][9] , \xmem_inst/mem[13][8] ,
         \xmem_inst/mem[13][7] , \xmem_inst/mem[13][6] ,
         \xmem_inst/mem[13][5] , \xmem_inst/mem[13][4] ,
         \xmem_inst/mem[13][3] , \xmem_inst/mem[13][2] ,
         \xmem_inst/mem[13][1] , \xmem_inst/mem[13][0] ,
         \xmem_inst/mem[12][31] , \xmem_inst/mem[12][30] ,
         \xmem_inst/mem[12][29] , \xmem_inst/mem[12][28] ,
         \xmem_inst/mem[12][27] , \xmem_inst/mem[12][26] ,
         \xmem_inst/mem[12][25] , \xmem_inst/mem[12][24] ,
         \xmem_inst/mem[12][23] , \xmem_inst/mem[12][22] ,
         \xmem_inst/mem[12][21] , \xmem_inst/mem[12][20] ,
         \xmem_inst/mem[12][19] , \xmem_inst/mem[12][18] ,
         \xmem_inst/mem[12][17] , \xmem_inst/mem[12][16] ,
         \xmem_inst/mem[12][15] , \xmem_inst/mem[12][14] ,
         \xmem_inst/mem[12][13] , \xmem_inst/mem[12][12] ,
         \xmem_inst/mem[12][11] , \xmem_inst/mem[12][10] ,
         \xmem_inst/mem[12][9] , \xmem_inst/mem[12][8] ,
         \xmem_inst/mem[12][7] , \xmem_inst/mem[12][6] ,
         \xmem_inst/mem[12][5] , \xmem_inst/mem[12][4] ,
         \xmem_inst/mem[12][3] , \xmem_inst/mem[12][2] ,
         \xmem_inst/mem[12][1] , \xmem_inst/mem[12][0] ,
         \xmem_inst/mem[11][31] , \xmem_inst/mem[11][30] ,
         \xmem_inst/mem[11][29] , \xmem_inst/mem[11][28] ,
         \xmem_inst/mem[11][27] , \xmem_inst/mem[11][26] ,
         \xmem_inst/mem[11][25] , \xmem_inst/mem[11][24] ,
         \xmem_inst/mem[11][23] , \xmem_inst/mem[11][22] ,
         \xmem_inst/mem[11][21] , \xmem_inst/mem[11][20] ,
         \xmem_inst/mem[11][19] , \xmem_inst/mem[11][18] ,
         \xmem_inst/mem[11][17] , \xmem_inst/mem[11][16] ,
         \xmem_inst/mem[11][15] , \xmem_inst/mem[11][14] ,
         \xmem_inst/mem[11][13] , \xmem_inst/mem[11][12] ,
         \xmem_inst/mem[11][11] , \xmem_inst/mem[11][10] ,
         \xmem_inst/mem[11][9] , \xmem_inst/mem[11][8] ,
         \xmem_inst/mem[11][7] , \xmem_inst/mem[11][6] ,
         \xmem_inst/mem[11][5] , \xmem_inst/mem[11][4] ,
         \xmem_inst/mem[11][3] , \xmem_inst/mem[11][2] ,
         \xmem_inst/mem[11][1] , \xmem_inst/mem[11][0] ,
         \xmem_inst/mem[10][31] , \xmem_inst/mem[10][30] ,
         \xmem_inst/mem[10][29] , \xmem_inst/mem[10][28] ,
         \xmem_inst/mem[10][27] , \xmem_inst/mem[10][26] ,
         \xmem_inst/mem[10][25] , \xmem_inst/mem[10][24] ,
         \xmem_inst/mem[10][23] , \xmem_inst/mem[10][22] ,
         \xmem_inst/mem[10][21] , \xmem_inst/mem[10][20] ,
         \xmem_inst/mem[10][19] , \xmem_inst/mem[10][18] ,
         \xmem_inst/mem[10][17] , \xmem_inst/mem[10][16] ,
         \xmem_inst/mem[10][15] , \xmem_inst/mem[10][14] ,
         \xmem_inst/mem[10][13] , \xmem_inst/mem[10][12] ,
         \xmem_inst/mem[10][11] , \xmem_inst/mem[10][10] ,
         \xmem_inst/mem[10][9] , \xmem_inst/mem[10][8] ,
         \xmem_inst/mem[10][7] , \xmem_inst/mem[10][6] ,
         \xmem_inst/mem[10][5] , \xmem_inst/mem[10][4] ,
         \xmem_inst/mem[10][3] , \xmem_inst/mem[10][2] ,
         \xmem_inst/mem[10][1] , \xmem_inst/mem[10][0] ,
         \xmem_inst/mem[9][31] , \xmem_inst/mem[9][30] ,
         \xmem_inst/mem[9][29] , \xmem_inst/mem[9][28] ,
         \xmem_inst/mem[9][27] , \xmem_inst/mem[9][26] ,
         \xmem_inst/mem[9][25] , \xmem_inst/mem[9][24] ,
         \xmem_inst/mem[9][23] , \xmem_inst/mem[9][22] ,
         \xmem_inst/mem[9][21] , \xmem_inst/mem[9][20] ,
         \xmem_inst/mem[9][19] , \xmem_inst/mem[9][18] ,
         \xmem_inst/mem[9][17] , \xmem_inst/mem[9][16] ,
         \xmem_inst/mem[9][15] , \xmem_inst/mem[9][14] ,
         \xmem_inst/mem[9][13] , \xmem_inst/mem[9][12] ,
         \xmem_inst/mem[9][11] , \xmem_inst/mem[9][10] , \xmem_inst/mem[9][9] ,
         \xmem_inst/mem[9][8] , \xmem_inst/mem[9][7] , \xmem_inst/mem[9][6] ,
         \xmem_inst/mem[9][5] , \xmem_inst/mem[9][4] , \xmem_inst/mem[9][3] ,
         \xmem_inst/mem[9][2] , \xmem_inst/mem[9][1] , \xmem_inst/mem[9][0] ,
         \xmem_inst/mem[8][31] , \xmem_inst/mem[8][30] ,
         \xmem_inst/mem[8][29] , \xmem_inst/mem[8][28] ,
         \xmem_inst/mem[8][27] , \xmem_inst/mem[8][26] ,
         \xmem_inst/mem[8][25] , \xmem_inst/mem[8][24] ,
         \xmem_inst/mem[8][23] , \xmem_inst/mem[8][22] ,
         \xmem_inst/mem[8][21] , \xmem_inst/mem[8][20] ,
         \xmem_inst/mem[8][19] , \xmem_inst/mem[8][18] ,
         \xmem_inst/mem[8][17] , \xmem_inst/mem[8][16] ,
         \xmem_inst/mem[8][15] , \xmem_inst/mem[8][14] ,
         \xmem_inst/mem[8][13] , \xmem_inst/mem[8][12] ,
         \xmem_inst/mem[8][11] , \xmem_inst/mem[8][10] , \xmem_inst/mem[8][9] ,
         \xmem_inst/mem[8][8] , \xmem_inst/mem[8][7] , \xmem_inst/mem[8][6] ,
         \xmem_inst/mem[8][5] , \xmem_inst/mem[8][4] , \xmem_inst/mem[8][3] ,
         \xmem_inst/mem[8][2] , \xmem_inst/mem[8][1] , \xmem_inst/mem[8][0] ,
         \xmem_inst/mem[7][31] , \xmem_inst/mem[7][30] ,
         \xmem_inst/mem[7][29] , \xmem_inst/mem[7][28] ,
         \xmem_inst/mem[7][27] , \xmem_inst/mem[7][26] ,
         \xmem_inst/mem[7][25] , \xmem_inst/mem[7][24] ,
         \xmem_inst/mem[7][23] , \xmem_inst/mem[7][22] ,
         \xmem_inst/mem[7][21] , \xmem_inst/mem[7][20] ,
         \xmem_inst/mem[7][19] , \xmem_inst/mem[7][18] ,
         \xmem_inst/mem[7][17] , \xmem_inst/mem[7][16] ,
         \xmem_inst/mem[7][15] , \xmem_inst/mem[7][14] ,
         \xmem_inst/mem[7][13] , \xmem_inst/mem[7][12] ,
         \xmem_inst/mem[7][11] , \xmem_inst/mem[7][10] , \xmem_inst/mem[7][9] ,
         \xmem_inst/mem[7][8] , \xmem_inst/mem[7][7] , \xmem_inst/mem[7][6] ,
         \xmem_inst/mem[7][5] , \xmem_inst/mem[7][4] , \xmem_inst/mem[7][3] ,
         \xmem_inst/mem[7][2] , \xmem_inst/mem[7][1] , \xmem_inst/mem[7][0] ,
         \xmem_inst/mem[6][31] , \xmem_inst/mem[6][30] ,
         \xmem_inst/mem[6][29] , \xmem_inst/mem[6][28] ,
         \xmem_inst/mem[6][27] , \xmem_inst/mem[6][26] ,
         \xmem_inst/mem[6][25] , \xmem_inst/mem[6][24] ,
         \xmem_inst/mem[6][23] , \xmem_inst/mem[6][22] ,
         \xmem_inst/mem[6][21] , \xmem_inst/mem[6][20] ,
         \xmem_inst/mem[6][19] , \xmem_inst/mem[6][18] ,
         \xmem_inst/mem[6][17] , \xmem_inst/mem[6][16] ,
         \xmem_inst/mem[6][15] , \xmem_inst/mem[6][14] ,
         \xmem_inst/mem[6][13] , \xmem_inst/mem[6][12] ,
         \xmem_inst/mem[6][11] , \xmem_inst/mem[6][10] , \xmem_inst/mem[6][9] ,
         \xmem_inst/mem[6][8] , \xmem_inst/mem[6][7] , \xmem_inst/mem[6][6] ,
         \xmem_inst/mem[6][5] , \xmem_inst/mem[6][4] , \xmem_inst/mem[6][3] ,
         \xmem_inst/mem[6][2] , \xmem_inst/mem[6][1] , \xmem_inst/mem[6][0] ,
         \xmem_inst/mem[5][31] , \xmem_inst/mem[5][30] ,
         \xmem_inst/mem[5][29] , \xmem_inst/mem[5][28] ,
         \xmem_inst/mem[5][27] , \xmem_inst/mem[5][26] ,
         \xmem_inst/mem[5][25] , \xmem_inst/mem[5][24] ,
         \xmem_inst/mem[5][23] , \xmem_inst/mem[5][22] ,
         \xmem_inst/mem[5][21] , \xmem_inst/mem[5][20] ,
         \xmem_inst/mem[5][19] , \xmem_inst/mem[5][18] ,
         \xmem_inst/mem[5][17] , \xmem_inst/mem[5][16] ,
         \xmem_inst/mem[5][15] , \xmem_inst/mem[5][14] ,
         \xmem_inst/mem[5][13] , \xmem_inst/mem[5][12] ,
         \xmem_inst/mem[5][11] , \xmem_inst/mem[5][10] , \xmem_inst/mem[5][9] ,
         \xmem_inst/mem[5][8] , \xmem_inst/mem[5][7] , \xmem_inst/mem[5][6] ,
         \xmem_inst/mem[5][5] , \xmem_inst/mem[5][4] , \xmem_inst/mem[5][3] ,
         \xmem_inst/mem[5][2] , \xmem_inst/mem[5][1] , \xmem_inst/mem[5][0] ,
         \xmem_inst/mem[4][31] , \xmem_inst/mem[4][30] ,
         \xmem_inst/mem[4][29] , \xmem_inst/mem[4][28] ,
         \xmem_inst/mem[4][27] , \xmem_inst/mem[4][26] ,
         \xmem_inst/mem[4][25] , \xmem_inst/mem[4][24] ,
         \xmem_inst/mem[4][23] , \xmem_inst/mem[4][22] ,
         \xmem_inst/mem[4][21] , \xmem_inst/mem[4][20] ,
         \xmem_inst/mem[4][19] , \xmem_inst/mem[4][18] ,
         \xmem_inst/mem[4][17] , \xmem_inst/mem[4][16] ,
         \xmem_inst/mem[4][15] , \xmem_inst/mem[4][14] ,
         \xmem_inst/mem[4][13] , \xmem_inst/mem[4][12] ,
         \xmem_inst/mem[4][11] , \xmem_inst/mem[4][10] , \xmem_inst/mem[4][9] ,
         \xmem_inst/mem[4][8] , \xmem_inst/mem[4][7] , \xmem_inst/mem[4][6] ,
         \xmem_inst/mem[4][5] , \xmem_inst/mem[4][4] , \xmem_inst/mem[4][3] ,
         \xmem_inst/mem[4][2] , \xmem_inst/mem[4][1] , \xmem_inst/mem[4][0] ,
         \xmem_inst/mem[3][31] , \xmem_inst/mem[3][30] ,
         \xmem_inst/mem[3][29] , \xmem_inst/mem[3][28] ,
         \xmem_inst/mem[3][27] , \xmem_inst/mem[3][26] ,
         \xmem_inst/mem[3][25] , \xmem_inst/mem[3][24] ,
         \xmem_inst/mem[3][23] , \xmem_inst/mem[3][22] ,
         \xmem_inst/mem[3][21] , \xmem_inst/mem[3][20] ,
         \xmem_inst/mem[3][19] , \xmem_inst/mem[3][18] ,
         \xmem_inst/mem[3][17] , \xmem_inst/mem[3][16] ,
         \xmem_inst/mem[3][15] , \xmem_inst/mem[3][14] ,
         \xmem_inst/mem[3][13] , \xmem_inst/mem[3][12] ,
         \xmem_inst/mem[3][11] , \xmem_inst/mem[3][10] , \xmem_inst/mem[3][9] ,
         \xmem_inst/mem[3][8] , \xmem_inst/mem[3][7] , \xmem_inst/mem[3][6] ,
         \xmem_inst/mem[3][5] , \xmem_inst/mem[3][4] , \xmem_inst/mem[3][3] ,
         \xmem_inst/mem[3][2] , \xmem_inst/mem[3][1] , \xmem_inst/mem[3][0] ,
         \xmem_inst/mem[2][31] , \xmem_inst/mem[2][30] ,
         \xmem_inst/mem[2][29] , \xmem_inst/mem[2][28] ,
         \xmem_inst/mem[2][27] , \xmem_inst/mem[2][26] ,
         \xmem_inst/mem[2][25] , \xmem_inst/mem[2][24] ,
         \xmem_inst/mem[2][23] , \xmem_inst/mem[2][22] ,
         \xmem_inst/mem[2][21] , \xmem_inst/mem[2][20] ,
         \xmem_inst/mem[2][19] , \xmem_inst/mem[2][18] ,
         \xmem_inst/mem[2][17] , \xmem_inst/mem[2][16] ,
         \xmem_inst/mem[2][15] , \xmem_inst/mem[2][14] ,
         \xmem_inst/mem[2][13] , \xmem_inst/mem[2][12] ,
         \xmem_inst/mem[2][11] , \xmem_inst/mem[2][10] , \xmem_inst/mem[2][9] ,
         \xmem_inst/mem[2][8] , \xmem_inst/mem[2][7] , \xmem_inst/mem[2][6] ,
         \xmem_inst/mem[2][5] , \xmem_inst/mem[2][4] , \xmem_inst/mem[2][3] ,
         \xmem_inst/mem[2][2] , \xmem_inst/mem[2][1] , \xmem_inst/mem[2][0] ,
         \xmem_inst/mem[1][31] , \xmem_inst/mem[1][30] ,
         \xmem_inst/mem[1][29] , \xmem_inst/mem[1][28] ,
         \xmem_inst/mem[1][27] , \xmem_inst/mem[1][26] ,
         \xmem_inst/mem[1][25] , \xmem_inst/mem[1][24] ,
         \xmem_inst/mem[1][23] , \xmem_inst/mem[1][22] ,
         \xmem_inst/mem[1][21] , \xmem_inst/mem[1][20] ,
         \xmem_inst/mem[1][19] , \xmem_inst/mem[1][18] ,
         \xmem_inst/mem[1][17] , \xmem_inst/mem[1][16] ,
         \xmem_inst/mem[1][15] , \xmem_inst/mem[1][14] ,
         \xmem_inst/mem[1][13] , \xmem_inst/mem[1][12] ,
         \xmem_inst/mem[1][11] , \xmem_inst/mem[1][10] , \xmem_inst/mem[1][9] ,
         \xmem_inst/mem[1][8] , \xmem_inst/mem[1][7] , \xmem_inst/mem[1][6] ,
         \xmem_inst/mem[1][5] , \xmem_inst/mem[1][4] , \xmem_inst/mem[1][3] ,
         \xmem_inst/mem[1][2] , \xmem_inst/mem[1][1] , \xmem_inst/mem[1][0] ,
         \xmem_inst/mem[0][31] , \xmem_inst/mem[0][30] ,
         \xmem_inst/mem[0][29] , \xmem_inst/mem[0][28] ,
         \xmem_inst/mem[0][27] , \xmem_inst/mem[0][26] ,
         \xmem_inst/mem[0][25] , \xmem_inst/mem[0][24] ,
         \xmem_inst/mem[0][23] , \xmem_inst/mem[0][22] ,
         \xmem_inst/mem[0][21] , \xmem_inst/mem[0][20] ,
         \xmem_inst/mem[0][19] , \xmem_inst/mem[0][18] ,
         \xmem_inst/mem[0][17] , \xmem_inst/mem[0][16] ,
         \xmem_inst/mem[0][15] , \xmem_inst/mem[0][14] ,
         \xmem_inst/mem[0][13] , \xmem_inst/mem[0][12] ,
         \xmem_inst/mem[0][11] , \xmem_inst/mem[0][10] , \xmem_inst/mem[0][9] ,
         \xmem_inst/mem[0][8] , \xmem_inst/mem[0][7] , \xmem_inst/mem[0][6] ,
         \xmem_inst/mem[0][5] , \xmem_inst/mem[0][4] , \xmem_inst/mem[0][3] ,
         \xmem_inst/mem[0][2] , \xmem_inst/mem[0][1] , \xmem_inst/mem[0][0] ,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2099, n2100, n2101, n2102, n2103, n2104, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362;
  wire   [5:0] xmem_addr;
  wire   [31:0] xmem_data;
  wire   [3:0] fmem_addr;
  wire   [31:0] fmem_data;
  wire   [5:0] \ctrl_conv_output_inst/cnt_conv ;
  wire   [31:0] \mac_unit_inst/adder_reg ;
  wire   [31:0] \mac_unit_inst/x_mult_f_reg ;
  assign m_data_out_y[31] = 1'b0;

  DFF_X1 \ctrl_conv_output_inst/conv_done_reg  ( .D(
        \ctrl_conv_output_inst/N80 ), .CK(clk), .Q(conv_done) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[5]  ( .D(n107), .CK(clk), .Q(
        xmem_addr[5]) );
  DFF_X1 conv_pre_start_reg ( .D(N23), .CK(clk), .Q(conv_pre_start) );
  DFF_X1 \ctrl_conv_output_inst/conv_start_accum_reg  ( .D(
        \ctrl_conv_output_inst/N77 ), .CK(clk), .Q(
        \ctrl_conv_output_inst/conv_start_accum ) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[0]  ( .D(\mac_unit_inst/n112 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [0]), .QN(n4084) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[1]  ( .D(\mac_unit_inst/n111 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [1]), .QN(n4085) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[2]  ( .D(\mac_unit_inst/n110 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [2]), .QN(n4086) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[3]  ( .D(\mac_unit_inst/n109 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [3]), .QN(n4087) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[4]  ( .D(\mac_unit_inst/n108 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [4]), .QN(n4103) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[5]  ( .D(\mac_unit_inst/n107 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [5]), .QN(n4104) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[6]  ( .D(\mac_unit_inst/n106 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [6]), .QN(n4088) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[7]  ( .D(\mac_unit_inst/n105 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [7]), .QN(n4089) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[8]  ( .D(\mac_unit_inst/n104 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [8]), .QN(n323) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[9]  ( .D(\mac_unit_inst/n103 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [9]), .QN(n324) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[10]  ( .D(\mac_unit_inst/n102 ), .CK(clk), .Q(\mac_unit_inst/adder_reg [10]), .QN(n322) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[11]  ( .D(\mac_unit_inst/n101 ), .CK(clk), .Q(\mac_unit_inst/adder_reg [11]), .QN(n325) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[12]  ( .D(\mac_unit_inst/n100 ), .CK(clk), .Q(\mac_unit_inst/adder_reg [12]), .QN(n4090) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[13]  ( .D(\mac_unit_inst/n99 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [13]), .QN(n4091) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[14]  ( .D(\mac_unit_inst/n98 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [14]), .QN(n4092) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[15]  ( .D(\mac_unit_inst/n97 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [15]), .QN(n4093) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[16]  ( .D(\mac_unit_inst/n96 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [16]), .QN(n4094) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[17]  ( .D(\mac_unit_inst/n95 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [17]), .QN(n4095) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[18]  ( .D(\mac_unit_inst/n94 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [18]), .QN(n4096) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[19]  ( .D(\mac_unit_inst/n93 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [19]), .QN(n4097) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[20]  ( .D(\mac_unit_inst/n92 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [20]), .QN(n4098) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[21]  ( .D(\mac_unit_inst/n91 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [21]), .QN(n4099) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[22]  ( .D(\mac_unit_inst/n90 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [22]), .QN(n4100) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[23]  ( .D(\mac_unit_inst/n89 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [23]), .QN(n4101) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[24]  ( .D(\mac_unit_inst/n88 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [24]), .QN(n326) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[25]  ( .D(\mac_unit_inst/n87 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [25]), .QN(n327) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[26]  ( .D(\mac_unit_inst/n86 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [26]), .QN(n328) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[27]  ( .D(\mac_unit_inst/n85 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [27]), .QN(n318) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[28]  ( .D(\mac_unit_inst/n84 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [28]), .QN(n319) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[29]  ( .D(\mac_unit_inst/n83 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [29]), .QN(n320) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[30]  ( .D(\mac_unit_inst/n82 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [30]), .QN(n321) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[0]  ( .D(\mac_unit_inst/n113 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [0]), .QN(n4144) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[1]  ( .D(\mac_unit_inst/n114 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [1]), .QN(n4119) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[2]  ( .D(\mac_unit_inst/n115 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [2]), .QN(n4118) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[3]  ( .D(\mac_unit_inst/n116 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [3]), .QN(n4117) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[4]  ( .D(\mac_unit_inst/n117 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [4]), .QN(n4116) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[5]  ( .D(\mac_unit_inst/n118 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [5]), .QN(n4115) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[6]  ( .D(\mac_unit_inst/n119 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [6]), .QN(n4114) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[7]  ( .D(\mac_unit_inst/n120 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [7]), .QN(n4131) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[8]  ( .D(\mac_unit_inst/n121 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [8]), .QN(n4130) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[9]  ( .D(\mac_unit_inst/n122 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [9]), .QN(n4129) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[10]  ( .D(\mac_unit_inst/n123 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [10]), .QN(n4128) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[11]  ( .D(\mac_unit_inst/n124 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [11]), .QN(n4127) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[12]  ( .D(\mac_unit_inst/n125 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [12]), .QN(n4126) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[13]  ( .D(\mac_unit_inst/n126 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [13]), .QN(n4125) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[14]  ( .D(\mac_unit_inst/n127 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [14]), .QN(n4124) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[15]  ( .D(\mac_unit_inst/n128 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [15]), .QN(n4123) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[16]  ( .D(\mac_unit_inst/n129 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [16]), .QN(n4122) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[17]  ( .D(\mac_unit_inst/n130 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [17]), .QN(n4121) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[18]  ( .D(\mac_unit_inst/n131 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [18]), .QN(n4120) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[20]  ( .D(\mac_unit_inst/n133 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [20]), .QN(n4142) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[21]  ( .D(\mac_unit_inst/n134 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [21]), .QN(n4141) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[22]  ( .D(\mac_unit_inst/n135 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [22]), .QN(n4140) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[25]  ( .D(\mac_unit_inst/n138 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [25]), .QN(n4137) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[26]  ( .D(\mac_unit_inst/n139 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [26]), .QN(n4136) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[27]  ( .D(\mac_unit_inst/n140 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [27]), .QN(n4135) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[28]  ( .D(\mac_unit_inst/n141 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [28]), .QN(n4134) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[29]  ( .D(\mac_unit_inst/n142 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [29]), .QN(n4133) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[30]  ( .D(\mac_unit_inst/n143 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [30]), .QN(n4132) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[31]  ( .D(\mac_unit_inst/n144 ), .CK(
        clk), .QN(n4112) );
  DFF_X1 \xmem_inst/data_out_reg[2]  ( .D(\xmem_inst/N277 ), .CK(clk), .Q(
        xmem_data[2]), .QN(n212) );
  DFF_X1 \xmem_inst/data_out_reg[4]  ( .D(\xmem_inst/N275 ), .CK(clk), .Q(
        xmem_data[4]) );
  DFF_X1 \xmem_inst/data_out_reg[5]  ( .D(\xmem_inst/N274 ), .CK(clk), .Q(
        xmem_data[5]), .QN(n4055) );
  DFF_X1 \xmem_inst/data_out_reg[6]  ( .D(\xmem_inst/N273 ), .CK(clk), .Q(n266), .QN(n4067) );
  DFF_X1 \xmem_inst/data_out_reg[7]  ( .D(\xmem_inst/N272 ), .CK(clk), .Q(
        xmem_data[7]), .QN(n4068) );
  DFF_X1 \xmem_inst/data_out_reg[8]  ( .D(\xmem_inst/N271 ), .CK(clk), .Q(
        xmem_data[8]), .QN(n270) );
  DFF_X1 \xmem_inst/data_out_reg[9]  ( .D(\xmem_inst/N270 ), .CK(clk), .Q(
        xmem_data[9]), .QN(n4051) );
  DFF_X1 \xmem_inst/data_out_reg[10]  ( .D(\xmem_inst/N269 ), .CK(clk), .Q(
        xmem_data[10]), .QN(n4050) );
  DFF_X1 \xmem_inst/data_out_reg[11]  ( .D(\xmem_inst/N268 ), .CK(clk), .Q(
        xmem_data[11]), .QN(n4058) );
  DFF_X1 \xmem_inst/data_out_reg[12]  ( .D(\xmem_inst/N267 ), .CK(clk), .Q(
        xmem_data[12]), .QN(n223) );
  DFF_X1 \xmem_inst/data_out_reg[13]  ( .D(\xmem_inst/N266 ), .CK(clk), .Q(
        xmem_data[13]), .QN(n4061) );
  DFF_X1 \xmem_inst/data_out_reg[14]  ( .D(\xmem_inst/N265 ), .CK(clk), .Q(
        xmem_data[14]), .QN(n333) );
  DFF_X1 \xmem_inst/data_out_reg[15]  ( .D(\xmem_inst/N264 ), .CK(clk), .Q(
        xmem_data[15]), .QN(n4053) );
  DFF_X1 \xmem_inst/data_out_reg[16]  ( .D(\xmem_inst/N263 ), .CK(clk), .QN(
        n269) );
  DFF_X1 \xmem_inst/data_out_reg[17]  ( .D(\xmem_inst/N262 ), .CK(clk), .Q(
        xmem_data[17]), .QN(n4059) );
  DFF_X1 \xmem_inst/data_out_reg[18]  ( .D(\xmem_inst/N261 ), .CK(clk), .Q(
        xmem_data[18]), .QN(n4060) );
  DFF_X1 \xmem_inst/data_out_reg[19]  ( .D(\xmem_inst/N260 ), .CK(clk), .Q(
        xmem_data[19]), .QN(n4064) );
  DFF_X1 \xmem_inst/data_out_reg[20]  ( .D(\xmem_inst/N259 ), .CK(clk), .QN(
        n4052) );
  DFF_X1 \xmem_inst/data_out_reg[22]  ( .D(\xmem_inst/N257 ), .CK(clk), .Q(
        xmem_data[22]), .QN(n221) );
  DFF_X1 \xmem_inst/data_out_reg[23]  ( .D(\xmem_inst/N256 ), .CK(clk), .Q(
        xmem_data[23]), .QN(n4062) );
  DFF_X1 \xmem_inst/data_out_reg[24]  ( .D(\xmem_inst/N255 ), .CK(clk), .QN(
        n313) );
  DFF_X1 \xmem_inst/data_out_reg[26]  ( .D(\xmem_inst/N253 ), .CK(clk), .Q(
        xmem_data[26]), .QN(n4066) );
  DFF_X1 \xmem_inst/data_out_reg[28]  ( .D(\xmem_inst/N251 ), .CK(clk), .Q(
        xmem_data[28]), .QN(n272) );
  DFF_X1 \xmem_inst/data_out_reg[30]  ( .D(\xmem_inst/N249 ), .CK(clk), .Q(
        xmem_data[30]) );
  DFF_X1 \xmem_inst/mem_reg[7][20]  ( .D(\xmem_inst/n2686 ), .CK(clk), .Q(
        \xmem_inst/mem[7][20] ), .QN(n4106) );
  DFF_X1 \xmem_inst/mem_reg[32][0]  ( .D(\xmem_inst/n3466 ), .CK(clk), .Q(
        \xmem_inst/mem[32][0] ) );
  DFF_X1 \xmem_inst/mem_reg[32][1]  ( .D(\xmem_inst/n3467 ), .CK(clk), .Q(
        \xmem_inst/mem[32][1] ) );
  DFF_X1 \xmem_inst/mem_reg[32][2]  ( .D(\xmem_inst/n3468 ), .CK(clk), .Q(
        \xmem_inst/mem[32][2] ) );
  DFF_X1 \xmem_inst/mem_reg[32][3]  ( .D(\xmem_inst/n3469 ), .CK(clk), .Q(
        \xmem_inst/mem[32][3] ) );
  DFF_X1 \xmem_inst/mem_reg[32][4]  ( .D(\xmem_inst/n3470 ), .CK(clk), .Q(
        \xmem_inst/mem[32][4] ) );
  DFF_X1 \xmem_inst/mem_reg[32][5]  ( .D(\xmem_inst/n3471 ), .CK(clk), .Q(
        \xmem_inst/mem[32][5] ) );
  DFF_X1 \xmem_inst/mem_reg[32][6]  ( .D(\xmem_inst/n3472 ), .CK(clk), .Q(
        \xmem_inst/mem[32][6] ) );
  DFF_X1 \xmem_inst/mem_reg[32][7]  ( .D(\xmem_inst/n3473 ), .CK(clk), .Q(
        \xmem_inst/mem[32][7] ) );
  DFF_X1 \xmem_inst/mem_reg[32][8]  ( .D(\xmem_inst/n3474 ), .CK(clk), .Q(
        \xmem_inst/mem[32][8] ) );
  DFF_X1 \xmem_inst/mem_reg[32][9]  ( .D(\xmem_inst/n3475 ), .CK(clk), .Q(
        \xmem_inst/mem[32][9] ) );
  DFF_X1 \xmem_inst/mem_reg[32][10]  ( .D(\xmem_inst/n3476 ), .CK(clk), .Q(
        \xmem_inst/mem[32][10] ) );
  DFF_X1 \xmem_inst/mem_reg[32][11]  ( .D(\xmem_inst/n3477 ), .CK(clk), .Q(
        \xmem_inst/mem[32][11] ) );
  DFF_X1 \xmem_inst/mem_reg[32][12]  ( .D(\xmem_inst/n3478 ), .CK(clk), .Q(
        \xmem_inst/mem[32][12] ) );
  DFF_X1 \xmem_inst/mem_reg[32][13]  ( .D(\xmem_inst/n3479 ), .CK(clk), .Q(
        \xmem_inst/mem[32][13] ) );
  DFF_X1 \xmem_inst/mem_reg[32][14]  ( .D(\xmem_inst/n3480 ), .CK(clk), .Q(
        \xmem_inst/mem[32][14] ) );
  DFF_X1 \xmem_inst/mem_reg[32][16]  ( .D(\xmem_inst/n3482 ), .CK(clk), .Q(
        \xmem_inst/mem[32][16] ) );
  DFF_X1 \xmem_inst/mem_reg[32][17]  ( .D(\xmem_inst/n3483 ), .CK(clk), .Q(
        \xmem_inst/mem[32][17] ) );
  DFF_X1 \xmem_inst/mem_reg[32][18]  ( .D(\xmem_inst/n3484 ), .CK(clk), .Q(
        \xmem_inst/mem[32][18] ) );
  DFF_X1 \xmem_inst/mem_reg[32][20]  ( .D(\xmem_inst/n3486 ), .CK(clk), .Q(
        \xmem_inst/mem[32][20] ) );
  DFF_X1 \xmem_inst/mem_reg[32][21]  ( .D(\xmem_inst/n3487 ), .CK(clk), .Q(
        \xmem_inst/mem[32][21] ) );
  DFF_X1 \xmem_inst/mem_reg[32][22]  ( .D(\xmem_inst/n3488 ), .CK(clk), .Q(
        \xmem_inst/mem[32][22] ) );
  DFF_X1 \xmem_inst/mem_reg[32][23]  ( .D(\xmem_inst/n3489 ), .CK(clk), .Q(
        \xmem_inst/mem[32][23] ) );
  DFF_X1 \xmem_inst/mem_reg[32][24]  ( .D(\xmem_inst/n3490 ), .CK(clk), .Q(
        \xmem_inst/mem[32][24] ) );
  DFF_X1 \xmem_inst/mem_reg[32][25]  ( .D(\xmem_inst/n3491 ), .CK(clk), .Q(
        \xmem_inst/mem[32][25] ) );
  DFF_X1 \xmem_inst/mem_reg[32][26]  ( .D(\xmem_inst/n3492 ), .CK(clk), .Q(
        \xmem_inst/mem[32][26] ) );
  DFF_X1 \xmem_inst/mem_reg[32][27]  ( .D(\xmem_inst/n3493 ), .CK(clk), .Q(
        \xmem_inst/mem[32][27] ) );
  DFF_X1 \xmem_inst/mem_reg[32][28]  ( .D(\xmem_inst/n3494 ), .CK(clk), .Q(
        \xmem_inst/mem[32][28] ) );
  DFF_X1 \xmem_inst/mem_reg[32][29]  ( .D(\xmem_inst/n3495 ), .CK(clk), .Q(
        \xmem_inst/mem[32][29] ) );
  DFF_X1 \xmem_inst/mem_reg[33][0]  ( .D(\xmem_inst/n3498 ), .CK(clk), .Q(
        \xmem_inst/mem[33][0] ) );
  DFF_X1 \xmem_inst/mem_reg[33][1]  ( .D(\xmem_inst/n3499 ), .CK(clk), .Q(
        \xmem_inst/mem[33][1] ) );
  DFF_X1 \xmem_inst/mem_reg[33][2]  ( .D(\xmem_inst/n3500 ), .CK(clk), .Q(
        \xmem_inst/mem[33][2] ) );
  DFF_X1 \xmem_inst/mem_reg[33][3]  ( .D(\xmem_inst/n3501 ), .CK(clk), .Q(
        \xmem_inst/mem[33][3] ) );
  DFF_X1 \xmem_inst/mem_reg[33][4]  ( .D(\xmem_inst/n3502 ), .CK(clk), .Q(
        \xmem_inst/mem[33][4] ) );
  DFF_X1 \xmem_inst/mem_reg[33][5]  ( .D(\xmem_inst/n3503 ), .CK(clk), .Q(
        \xmem_inst/mem[33][5] ) );
  DFF_X1 \xmem_inst/mem_reg[33][6]  ( .D(\xmem_inst/n3504 ), .CK(clk), .Q(
        \xmem_inst/mem[33][6] ) );
  DFF_X1 \xmem_inst/mem_reg[33][7]  ( .D(\xmem_inst/n3505 ), .CK(clk), .Q(
        \xmem_inst/mem[33][7] ) );
  DFF_X1 \xmem_inst/mem_reg[33][8]  ( .D(\xmem_inst/n3506 ), .CK(clk), .Q(
        \xmem_inst/mem[33][8] ) );
  DFF_X1 \xmem_inst/mem_reg[33][9]  ( .D(\xmem_inst/n3507 ), .CK(clk), .Q(
        \xmem_inst/mem[33][9] ) );
  DFF_X1 \xmem_inst/mem_reg[33][10]  ( .D(\xmem_inst/n3508 ), .CK(clk), .Q(
        \xmem_inst/mem[33][10] ) );
  DFF_X1 \xmem_inst/mem_reg[33][11]  ( .D(\xmem_inst/n3509 ), .CK(clk), .Q(
        \xmem_inst/mem[33][11] ) );
  DFF_X1 \xmem_inst/mem_reg[33][12]  ( .D(\xmem_inst/n3510 ), .CK(clk), .Q(
        \xmem_inst/mem[33][12] ) );
  DFF_X1 \xmem_inst/mem_reg[33][13]  ( .D(\xmem_inst/n3511 ), .CK(clk), .Q(
        \xmem_inst/mem[33][13] ) );
  DFF_X1 \xmem_inst/mem_reg[33][14]  ( .D(\xmem_inst/n3512 ), .CK(clk), .Q(
        \xmem_inst/mem[33][14] ) );
  DFF_X1 \xmem_inst/mem_reg[33][16]  ( .D(\xmem_inst/n3514 ), .CK(clk), .Q(
        \xmem_inst/mem[33][16] ) );
  DFF_X1 \xmem_inst/mem_reg[33][17]  ( .D(\xmem_inst/n3515 ), .CK(clk), .Q(
        \xmem_inst/mem[33][17] ) );
  DFF_X1 \xmem_inst/mem_reg[33][18]  ( .D(\xmem_inst/n3516 ), .CK(clk), .Q(
        \xmem_inst/mem[33][18] ) );
  DFF_X1 \xmem_inst/mem_reg[33][25]  ( .D(\xmem_inst/n3523 ), .CK(clk), .Q(
        \xmem_inst/mem[33][25] ) );
  DFF_X1 \xmem_inst/mem_reg[33][27]  ( .D(\xmem_inst/n3525 ), .CK(clk), .Q(
        \xmem_inst/mem[33][27] ) );
  DFF_X1 \xmem_inst/mem_reg[33][29]  ( .D(\xmem_inst/n3527 ), .CK(clk), .Q(
        \xmem_inst/mem[33][29] ) );
  DFF_X1 \xmem_inst/mem_reg[34][5]  ( .D(\xmem_inst/n3535 ), .CK(clk), .Q(
        \xmem_inst/mem[34][5] ) );
  DFF_X1 \xmem_inst/mem_reg[34][6]  ( .D(\xmem_inst/n3536 ), .CK(clk), .Q(
        \xmem_inst/mem[34][6] ) );
  DFF_X1 \xmem_inst/mem_reg[34][7]  ( .D(\xmem_inst/n3537 ), .CK(clk), .Q(
        \xmem_inst/mem[34][7] ) );
  DFF_X1 \xmem_inst/mem_reg[34][8]  ( .D(\xmem_inst/n3538 ), .CK(clk), .Q(
        \xmem_inst/mem[34][8] ) );
  DFF_X1 \xmem_inst/mem_reg[34][9]  ( .D(\xmem_inst/n3539 ), .CK(clk), .Q(
        \xmem_inst/mem[34][9] ) );
  DFF_X1 \xmem_inst/mem_reg[34][11]  ( .D(\xmem_inst/n3541 ), .CK(clk), .Q(
        \xmem_inst/mem[34][11] ) );
  DFF_X1 \xmem_inst/mem_reg[34][14]  ( .D(\xmem_inst/n3544 ), .CK(clk), .Q(
        \xmem_inst/mem[34][14] ) );
  DFF_X1 \xmem_inst/mem_reg[34][25]  ( .D(\xmem_inst/n3555 ), .CK(clk), .Q(
        \xmem_inst/mem[34][25] ) );
  DFF_X1 \xmem_inst/mem_reg[34][27]  ( .D(\xmem_inst/n3557 ), .CK(clk), .Q(
        \xmem_inst/mem[34][27] ) );
  DFF_X1 \xmem_inst/mem_reg[34][29]  ( .D(\xmem_inst/n3559 ), .CK(clk), .Q(
        \xmem_inst/mem[34][29] ) );
  DFF_X1 \xmem_inst/mem_reg[35][12]  ( .D(\xmem_inst/n3574 ), .CK(clk), .Q(
        \xmem_inst/mem[35][12] ), .QN(n4107) );
  DFF_X1 \xmem_inst/mem_reg[39][4]  ( .D(\xmem_inst/n3694 ), .CK(clk), .Q(
        \xmem_inst/mem[39][4] ), .QN(n4109) );
  DFF_X1 \xmem_inst/mem_reg[40][0]  ( .D(\xmem_inst/n3722 ), .CK(clk), .Q(
        \xmem_inst/mem[40][0] ) );
  DFF_X1 \xmem_inst/mem_reg[40][1]  ( .D(\xmem_inst/n3723 ), .CK(clk), .Q(
        \xmem_inst/mem[40][1] ) );
  DFF_X1 \xmem_inst/mem_reg[40][2]  ( .D(\xmem_inst/n3724 ), .CK(clk), .Q(
        \xmem_inst/mem[40][2] ) );
  DFF_X1 \xmem_inst/mem_reg[40][3]  ( .D(\xmem_inst/n3725 ), .CK(clk), .Q(
        \xmem_inst/mem[40][3] ) );
  DFF_X1 \xmem_inst/mem_reg[40][4]  ( .D(\xmem_inst/n3726 ), .CK(clk), .Q(
        \xmem_inst/mem[40][4] ) );
  DFF_X1 \xmem_inst/mem_reg[40][5]  ( .D(\xmem_inst/n3727 ), .CK(clk), .Q(
        \xmem_inst/mem[40][5] ) );
  DFF_X1 \xmem_inst/mem_reg[40][6]  ( .D(\xmem_inst/n3728 ), .CK(clk), .Q(
        \xmem_inst/mem[40][6] ) );
  DFF_X1 \xmem_inst/mem_reg[40][7]  ( .D(\xmem_inst/n3729 ), .CK(clk), .Q(
        \xmem_inst/mem[40][7] ) );
  DFF_X1 \xmem_inst/mem_reg[40][8]  ( .D(\xmem_inst/n3730 ), .CK(clk), .Q(
        \xmem_inst/mem[40][8] ) );
  DFF_X1 \xmem_inst/mem_reg[40][9]  ( .D(\xmem_inst/n3731 ), .CK(clk), .Q(
        \xmem_inst/mem[40][9] ) );
  DFF_X1 \xmem_inst/mem_reg[40][10]  ( .D(\xmem_inst/n3732 ), .CK(clk), .Q(
        \xmem_inst/mem[40][10] ) );
  DFF_X1 \xmem_inst/mem_reg[40][11]  ( .D(\xmem_inst/n3733 ), .CK(clk), .Q(
        \xmem_inst/mem[40][11] ) );
  DFF_X1 \xmem_inst/mem_reg[40][12]  ( .D(\xmem_inst/n3734 ), .CK(clk), .Q(
        \xmem_inst/mem[40][12] ) );
  DFF_X1 \xmem_inst/mem_reg[40][13]  ( .D(\xmem_inst/n3735 ), .CK(clk), .Q(
        \xmem_inst/mem[40][13] ) );
  DFF_X1 \xmem_inst/mem_reg[40][14]  ( .D(\xmem_inst/n3736 ), .CK(clk), .Q(
        \xmem_inst/mem[40][14] ) );
  DFF_X1 \xmem_inst/mem_reg[40][15]  ( .D(\xmem_inst/n3737 ), .CK(clk), .Q(
        \xmem_inst/mem[40][15] ) );
  DFF_X1 \xmem_inst/mem_reg[40][16]  ( .D(\xmem_inst/n3738 ), .CK(clk), .Q(
        \xmem_inst/mem[40][16] ) );
  DFF_X1 \xmem_inst/mem_reg[40][17]  ( .D(\xmem_inst/n3739 ), .CK(clk), .Q(
        \xmem_inst/mem[40][17] ) );
  DFF_X1 \xmem_inst/mem_reg[40][18]  ( .D(\xmem_inst/n3740 ), .CK(clk), .Q(
        \xmem_inst/mem[40][18] ) );
  DFF_X1 \xmem_inst/mem_reg[40][19]  ( .D(\xmem_inst/n3741 ), .CK(clk), .Q(
        \xmem_inst/mem[40][19] ) );
  DFF_X1 \xmem_inst/mem_reg[40][20]  ( .D(\xmem_inst/n3742 ), .CK(clk), .Q(
        \xmem_inst/mem[40][20] ) );
  DFF_X1 \xmem_inst/mem_reg[40][21]  ( .D(\xmem_inst/n3743 ), .CK(clk), .Q(
        \xmem_inst/mem[40][21] ) );
  DFF_X1 \xmem_inst/mem_reg[40][22]  ( .D(\xmem_inst/n3744 ), .CK(clk), .Q(
        \xmem_inst/mem[40][22] ) );
  DFF_X1 \xmem_inst/mem_reg[40][23]  ( .D(\xmem_inst/n3745 ), .CK(clk), .Q(
        \xmem_inst/mem[40][23] ) );
  DFF_X1 \xmem_inst/mem_reg[40][24]  ( .D(\xmem_inst/n3746 ), .CK(clk), .Q(
        \xmem_inst/mem[40][24] ) );
  DFF_X1 \xmem_inst/mem_reg[40][25]  ( .D(\xmem_inst/n3747 ), .CK(clk), .Q(
        \xmem_inst/mem[40][25] ) );
  DFF_X1 \xmem_inst/mem_reg[40][26]  ( .D(\xmem_inst/n3748 ), .CK(clk), .Q(
        \xmem_inst/mem[40][26] ) );
  DFF_X1 \xmem_inst/mem_reg[40][27]  ( .D(\xmem_inst/n3749 ), .CK(clk), .Q(
        \xmem_inst/mem[40][27] ) );
  DFF_X1 \xmem_inst/mem_reg[40][28]  ( .D(\xmem_inst/n3750 ), .CK(clk), .Q(
        \xmem_inst/mem[40][28] ) );
  DFF_X1 \xmem_inst/mem_reg[40][29]  ( .D(\xmem_inst/n3751 ), .CK(clk), .Q(
        \xmem_inst/mem[40][29] ) );
  DFF_X1 \xmem_inst/mem_reg[40][30]  ( .D(\xmem_inst/n3752 ), .CK(clk), .Q(
        \xmem_inst/mem[40][30] ) );
  DFF_X1 \xmem_inst/mem_reg[40][31]  ( .D(\xmem_inst/n3753 ), .CK(clk), .Q(
        \xmem_inst/mem[40][31] ) );
  DFF_X1 \xmem_inst/mem_reg[41][0]  ( .D(\xmem_inst/n3754 ), .CK(clk), .Q(
        \xmem_inst/mem[41][0] ) );
  DFF_X1 \xmem_inst/mem_reg[41][1]  ( .D(\xmem_inst/n3755 ), .CK(clk), .Q(
        \xmem_inst/mem[41][1] ) );
  DFF_X1 \xmem_inst/mem_reg[41][2]  ( .D(\xmem_inst/n3756 ), .CK(clk), .Q(
        \xmem_inst/mem[41][2] ) );
  DFF_X1 \xmem_inst/mem_reg[41][3]  ( .D(\xmem_inst/n3757 ), .CK(clk), .Q(
        \xmem_inst/mem[41][3] ) );
  DFF_X1 \xmem_inst/mem_reg[41][4]  ( .D(\xmem_inst/n3758 ), .CK(clk), .Q(
        \xmem_inst/mem[41][4] ) );
  DFF_X1 \xmem_inst/mem_reg[41][5]  ( .D(\xmem_inst/n3759 ), .CK(clk), .Q(
        \xmem_inst/mem[41][5] ) );
  DFF_X1 \xmem_inst/mem_reg[41][6]  ( .D(\xmem_inst/n3760 ), .CK(clk), .Q(
        \xmem_inst/mem[41][6] ) );
  DFF_X1 \xmem_inst/mem_reg[41][7]  ( .D(\xmem_inst/n3761 ), .CK(clk), .Q(
        \xmem_inst/mem[41][7] ) );
  DFF_X1 \xmem_inst/mem_reg[41][8]  ( .D(\xmem_inst/n3762 ), .CK(clk), .Q(
        \xmem_inst/mem[41][8] ) );
  DFF_X1 \xmem_inst/mem_reg[41][9]  ( .D(\xmem_inst/n3763 ), .CK(clk), .Q(
        \xmem_inst/mem[41][9] ) );
  DFF_X1 \xmem_inst/mem_reg[41][10]  ( .D(\xmem_inst/n3764 ), .CK(clk), .Q(
        \xmem_inst/mem[41][10] ) );
  DFF_X1 \xmem_inst/mem_reg[41][11]  ( .D(\xmem_inst/n3765 ), .CK(clk), .Q(
        \xmem_inst/mem[41][11] ) );
  DFF_X1 \xmem_inst/mem_reg[41][12]  ( .D(\xmem_inst/n3766 ), .CK(clk), .Q(
        \xmem_inst/mem[41][12] ) );
  DFF_X1 \xmem_inst/mem_reg[41][13]  ( .D(\xmem_inst/n3767 ), .CK(clk), .Q(
        \xmem_inst/mem[41][13] ) );
  DFF_X1 \xmem_inst/mem_reg[41][14]  ( .D(\xmem_inst/n3768 ), .CK(clk), .Q(
        \xmem_inst/mem[41][14] ) );
  DFF_X1 \xmem_inst/mem_reg[41][15]  ( .D(\xmem_inst/n3769 ), .CK(clk), .Q(
        \xmem_inst/mem[41][15] ) );
  DFF_X1 \xmem_inst/mem_reg[41][16]  ( .D(\xmem_inst/n3770 ), .CK(clk), .Q(
        \xmem_inst/mem[41][16] ) );
  DFF_X1 \xmem_inst/mem_reg[41][17]  ( .D(\xmem_inst/n3771 ), .CK(clk), .Q(
        \xmem_inst/mem[41][17] ) );
  DFF_X1 \xmem_inst/mem_reg[41][18]  ( .D(\xmem_inst/n3772 ), .CK(clk), .Q(
        \xmem_inst/mem[41][18] ) );
  DFF_X1 \xmem_inst/mem_reg[41][19]  ( .D(\xmem_inst/n3773 ), .CK(clk), .Q(
        \xmem_inst/mem[41][19] ) );
  DFF_X1 \xmem_inst/mem_reg[41][20]  ( .D(\xmem_inst/n3774 ), .CK(clk), .Q(
        \xmem_inst/mem[41][20] ) );
  DFF_X1 \xmem_inst/mem_reg[41][21]  ( .D(\xmem_inst/n3775 ), .CK(clk), .Q(
        \xmem_inst/mem[41][21] ) );
  DFF_X1 \xmem_inst/mem_reg[41][22]  ( .D(\xmem_inst/n3776 ), .CK(clk), .Q(
        \xmem_inst/mem[41][22] ) );
  DFF_X1 \xmem_inst/mem_reg[41][23]  ( .D(\xmem_inst/n3777 ), .CK(clk), .Q(
        \xmem_inst/mem[41][23] ) );
  DFF_X1 \xmem_inst/mem_reg[41][24]  ( .D(\xmem_inst/n3778 ), .CK(clk), .Q(
        \xmem_inst/mem[41][24] ) );
  DFF_X1 \xmem_inst/mem_reg[41][25]  ( .D(\xmem_inst/n3779 ), .CK(clk), .Q(
        \xmem_inst/mem[41][25] ) );
  DFF_X1 \xmem_inst/mem_reg[41][26]  ( .D(\xmem_inst/n3780 ), .CK(clk), .Q(
        \xmem_inst/mem[41][26] ) );
  DFF_X1 \xmem_inst/mem_reg[41][27]  ( .D(\xmem_inst/n3781 ), .CK(clk), .Q(
        \xmem_inst/mem[41][27] ) );
  DFF_X1 \xmem_inst/mem_reg[41][28]  ( .D(\xmem_inst/n3782 ), .CK(clk), .Q(
        \xmem_inst/mem[41][28] ) );
  DFF_X1 \xmem_inst/mem_reg[41][29]  ( .D(\xmem_inst/n3783 ), .CK(clk), .Q(
        \xmem_inst/mem[41][29] ) );
  DFF_X1 \xmem_inst/mem_reg[41][30]  ( .D(\xmem_inst/n3784 ), .CK(clk), .Q(
        \xmem_inst/mem[41][30] ) );
  DFF_X1 \xmem_inst/mem_reg[41][31]  ( .D(\xmem_inst/n3785 ), .CK(clk), .Q(
        \xmem_inst/mem[41][31] ) );
  DFF_X1 \xmem_inst/mem_reg[42][0]  ( .D(\xmem_inst/n3786 ), .CK(clk), .Q(
        \xmem_inst/mem[42][0] ) );
  DFF_X1 \xmem_inst/mem_reg[42][1]  ( .D(\xmem_inst/n3787 ), .CK(clk), .Q(
        \xmem_inst/mem[42][1] ) );
  DFF_X1 \xmem_inst/mem_reg[42][2]  ( .D(\xmem_inst/n3788 ), .CK(clk), .Q(
        \xmem_inst/mem[42][2] ) );
  DFF_X1 \xmem_inst/mem_reg[42][3]  ( .D(\xmem_inst/n3789 ), .CK(clk), .Q(
        \xmem_inst/mem[42][3] ) );
  DFF_X1 \xmem_inst/mem_reg[42][4]  ( .D(\xmem_inst/n3790 ), .CK(clk), .Q(
        \xmem_inst/mem[42][4] ) );
  DFF_X1 \xmem_inst/mem_reg[42][5]  ( .D(\xmem_inst/n3791 ), .CK(clk), .Q(
        \xmem_inst/mem[42][5] ) );
  DFF_X1 \xmem_inst/mem_reg[42][6]  ( .D(\xmem_inst/n3792 ), .CK(clk), .Q(
        \xmem_inst/mem[42][6] ) );
  DFF_X1 \xmem_inst/mem_reg[42][7]  ( .D(\xmem_inst/n3793 ), .CK(clk), .Q(
        \xmem_inst/mem[42][7] ) );
  DFF_X1 \xmem_inst/mem_reg[42][8]  ( .D(\xmem_inst/n3794 ), .CK(clk), .Q(
        \xmem_inst/mem[42][8] ) );
  DFF_X1 \xmem_inst/mem_reg[42][9]  ( .D(\xmem_inst/n3795 ), .CK(clk), .Q(
        \xmem_inst/mem[42][9] ) );
  DFF_X1 \xmem_inst/mem_reg[42][10]  ( .D(\xmem_inst/n3796 ), .CK(clk), .Q(
        \xmem_inst/mem[42][10] ) );
  DFF_X1 \xmem_inst/mem_reg[42][11]  ( .D(\xmem_inst/n3797 ), .CK(clk), .Q(
        \xmem_inst/mem[42][11] ) );
  DFF_X1 \xmem_inst/mem_reg[42][12]  ( .D(\xmem_inst/n3798 ), .CK(clk), .Q(
        \xmem_inst/mem[42][12] ) );
  DFF_X1 \xmem_inst/mem_reg[42][13]  ( .D(\xmem_inst/n3799 ), .CK(clk), .Q(
        \xmem_inst/mem[42][13] ) );
  DFF_X1 \xmem_inst/mem_reg[42][14]  ( .D(\xmem_inst/n3800 ), .CK(clk), .Q(
        \xmem_inst/mem[42][14] ) );
  DFF_X1 \xmem_inst/mem_reg[42][15]  ( .D(\xmem_inst/n3801 ), .CK(clk), .Q(
        \xmem_inst/mem[42][15] ) );
  DFF_X1 \xmem_inst/mem_reg[42][16]  ( .D(\xmem_inst/n3802 ), .CK(clk), .Q(
        \xmem_inst/mem[42][16] ) );
  DFF_X1 \xmem_inst/mem_reg[42][17]  ( .D(\xmem_inst/n3803 ), .CK(clk), .Q(
        \xmem_inst/mem[42][17] ) );
  DFF_X1 \xmem_inst/mem_reg[42][18]  ( .D(\xmem_inst/n3804 ), .CK(clk), .Q(
        \xmem_inst/mem[42][18] ) );
  DFF_X1 \xmem_inst/mem_reg[42][19]  ( .D(\xmem_inst/n3805 ), .CK(clk), .Q(
        \xmem_inst/mem[42][19] ) );
  DFF_X1 \xmem_inst/mem_reg[42][20]  ( .D(\xmem_inst/n3806 ), .CK(clk), .Q(
        \xmem_inst/mem[42][20] ) );
  DFF_X1 \xmem_inst/mem_reg[42][21]  ( .D(\xmem_inst/n3807 ), .CK(clk), .Q(
        \xmem_inst/mem[42][21] ) );
  DFF_X1 \xmem_inst/mem_reg[42][22]  ( .D(\xmem_inst/n3808 ), .CK(clk), .Q(
        \xmem_inst/mem[42][22] ) );
  DFF_X1 \xmem_inst/mem_reg[42][23]  ( .D(\xmem_inst/n3809 ), .CK(clk), .Q(
        \xmem_inst/mem[42][23] ) );
  DFF_X1 \xmem_inst/mem_reg[42][24]  ( .D(\xmem_inst/n3810 ), .CK(clk), .Q(
        \xmem_inst/mem[42][24] ) );
  DFF_X1 \xmem_inst/mem_reg[42][25]  ( .D(\xmem_inst/n3811 ), .CK(clk), .Q(
        \xmem_inst/mem[42][25] ) );
  DFF_X1 \xmem_inst/mem_reg[42][26]  ( .D(\xmem_inst/n3812 ), .CK(clk), .Q(
        \xmem_inst/mem[42][26] ) );
  DFF_X1 \xmem_inst/mem_reg[42][27]  ( .D(\xmem_inst/n3813 ), .CK(clk), .Q(
        \xmem_inst/mem[42][27] ) );
  DFF_X1 \xmem_inst/mem_reg[42][28]  ( .D(\xmem_inst/n3814 ), .CK(clk), .Q(
        \xmem_inst/mem[42][28] ) );
  DFF_X1 \xmem_inst/mem_reg[42][29]  ( .D(\xmem_inst/n3815 ), .CK(clk), .Q(
        \xmem_inst/mem[42][29] ) );
  DFF_X1 \xmem_inst/mem_reg[42][30]  ( .D(\xmem_inst/n3816 ), .CK(clk), .Q(
        \xmem_inst/mem[42][30] ) );
  DFF_X1 \xmem_inst/mem_reg[42][31]  ( .D(\xmem_inst/n3817 ), .CK(clk), .Q(
        \xmem_inst/mem[42][31] ) );
  DFF_X1 \xmem_inst/data_out_reg[21]  ( .D(\xmem_inst/N258 ), .CK(clk), .Q(
        xmem_data[21]), .QN(n330) );
  DFF_X1 \xmem_inst/data_out_reg[1]  ( .D(\xmem_inst/N278 ), .CK(clk), .Q(
        xmem_data[1]), .QN(n339) );
  DFF_X1 \xmem_inst/data_out_reg[3]  ( .D(\xmem_inst/N276 ), .CK(clk), .Q(
        xmem_data[3]), .QN(n329) );
  DFF_X1 \xmem_inst/data_out_reg[27]  ( .D(\xmem_inst/N252 ), .CK(clk), .Q(
        xmem_data[27]), .QN(n312) );
  DFF_X2 \xmem_inst/data_out_reg[31]  ( .D(\xmem_inst/N248 ), .CK(clk), .Q(
        xmem_data[31]), .QN(n4054) );
  DFF_X1 \xmem_inst/data_out_reg[29]  ( .D(\xmem_inst/N250 ), .CK(clk), .Q(
        xmem_data[29]), .QN(n331) );
  DFF_X1 \fmem_inst/z_reg[31]  ( .D(\fmem_inst/N78 ), .CK(clk), .Q(
        fmem_data[31]) );
  DFF_X1 \xmem_inst/data_out_reg[25]  ( .D(\xmem_inst/N254 ), .CK(clk), .Q(
        xmem_data[25]), .QN(n4065) );
  DFF_X2 \fmem_inst/z_reg[9]  ( .D(\fmem_inst/N71 ), .CK(clk), .Q(fmem_data[9]), .QN(n4057) );
  DFF_X2 \fmem_inst/z_reg[12]  ( .D(\fmem_inst/N74 ), .CK(clk), .Q(
        fmem_data[12]), .QN(n4056) );
  DFF_X2 \fmem_inst/z_reg[8]  ( .D(\fmem_inst/N70 ), .CK(clk), .Q(fmem_data[8]), .QN(n257) );
  DFF_X2 \fmem_inst/z_reg[5]  ( .D(\fmem_inst/N67 ), .CK(clk), .Q(fmem_data[5]), .QN(n273) );
  DFF_X2 \fmem_inst/z_reg[11]  ( .D(\fmem_inst/N73 ), .CK(clk), .Q(
        fmem_data[11]), .QN(n271) );
  DFF_X1 \ctrl_conv_output_inst/m_pre_pre_valid_y_reg  ( .D(n121), .CK(clk), 
        .Q(\ctrl_conv_output_inst/m_pre_pre_valid_y ), .QN(n4071) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[0]  ( .D(n119), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [0]), .QN(n4072) );
  DFF_X1 \ctrl_conv_output_inst/m_pre_valid_y_reg  ( .D(n106), .CK(clk), .Q(
        \ctrl_conv_output_inst/m_pre_valid_y ), .QN(n4075) );
  DFF_X1 \ctrl_conv_output_inst/m_valid_y_reg  ( .D(n114), .CK(clk), .Q(
        m_valid_y), .QN(n4073) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[3]  ( .D(n116), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [3]), .QN(n4110) );
  DFF_X1 \ctrl_xmem_write_inst/s_ready_reg  ( .D(n113), .CK(clk), .Q(s_ready_x), .QN(n4102) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[2]  ( .D(n117), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [2]), .QN(n4080) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[1]  ( .D(n118), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [1]), .QN(n4079) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[4]  ( .D(n115), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [4]), .QN(n4076) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[5]  ( .D(n120), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [5]), .QN(n4111) );
  DFF_X1 \fmem_addr_reg[0]  ( .D(n104), .CK(clk), .Q(fmem_addr[0]), .QN(n4074)
         );
  DFF_X1 \fmem_addr_reg[2]  ( .D(n102), .CK(clk), .Q(fmem_addr[2]), .QN(n4078)
         );
  DFF_X1 \fmem_addr_reg[1]  ( .D(n103), .CK(clk), .Q(fmem_addr[1]), .QN(n4069)
         );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[0]  ( .D(n112), .CK(clk), .Q(
        xmem_addr[0]), .QN(n4082) );
  DFF_X1 \fmem_addr_reg[3]  ( .D(n105), .CK(clk), .Q(fmem_addr[3]), .QN(n4077)
         );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[1]  ( .D(n111), .CK(clk), .Q(
        xmem_addr[1]), .QN(n4070) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[3]  ( .D(n109), .CK(clk), .Q(
        xmem_addr[3]), .QN(n4083) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[4]  ( .D(n108), .CK(clk), .Q(
        xmem_addr[4]), .QN(n4081) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[2]  ( .D(n4113), .CK(clk), .Q(
        n4105), .QN(xmem_addr[2]) );
  DFF_X1 \xmem_inst/mem_reg[7][8]  ( .D(n4377), .CK(clk), .Q(n4108), .QN(
        \xmem_inst/mem[7][8] ) );
  DFF_X1 \xmem_inst/mem_reg[23][31]  ( .D(n4911), .CK(clk), .QN(
        \xmem_inst/mem[23][31] ) );
  DFF_X1 \xmem_inst/mem_reg[23][30]  ( .D(n4910), .CK(clk), .QN(
        \xmem_inst/mem[23][30] ) );
  DFF_X1 \xmem_inst/mem_reg[23][19]  ( .D(n4899), .CK(clk), .QN(
        \xmem_inst/mem[23][19] ) );
  DFF_X1 \xmem_inst/mem_reg[23][15]  ( .D(n4895), .CK(clk), .QN(
        \xmem_inst/mem[23][15] ) );
  DFF_X1 \xmem_inst/mem_reg[22][31]  ( .D(n4879), .CK(clk), .QN(
        \xmem_inst/mem[22][31] ) );
  DFF_X1 \xmem_inst/mem_reg[22][30]  ( .D(n4878), .CK(clk), .QN(
        \xmem_inst/mem[22][30] ) );
  DFF_X1 \xmem_inst/mem_reg[22][19]  ( .D(n4867), .CK(clk), .QN(
        \xmem_inst/mem[22][19] ) );
  DFF_X1 \xmem_inst/mem_reg[22][15]  ( .D(n4863), .CK(clk), .QN(
        \xmem_inst/mem[22][15] ) );
  DFF_X1 \xmem_inst/mem_reg[21][31]  ( .D(n4847), .CK(clk), .QN(
        \xmem_inst/mem[21][31] ) );
  DFF_X1 \xmem_inst/mem_reg[21][30]  ( .D(n4846), .CK(clk), .QN(
        \xmem_inst/mem[21][30] ) );
  DFF_X1 \xmem_inst/mem_reg[21][19]  ( .D(n4835), .CK(clk), .QN(
        \xmem_inst/mem[21][19] ) );
  DFF_X1 \xmem_inst/mem_reg[21][15]  ( .D(n4831), .CK(clk), .QN(
        \xmem_inst/mem[21][15] ) );
  DFF_X1 \xmem_inst/mem_reg[20][31]  ( .D(n4815), .CK(clk), .QN(
        \xmem_inst/mem[20][31] ) );
  DFF_X1 \xmem_inst/mem_reg[20][30]  ( .D(n4814), .CK(clk), .QN(
        \xmem_inst/mem[20][30] ) );
  DFF_X1 \xmem_inst/mem_reg[20][19]  ( .D(n4803), .CK(clk), .QN(
        \xmem_inst/mem[20][19] ) );
  DFF_X1 \xmem_inst/mem_reg[20][15]  ( .D(n4799), .CK(clk), .QN(
        \xmem_inst/mem[20][15] ) );
  DFF_X1 \xmem_inst/mem_reg[19][31]  ( .D(n4783), .CK(clk), .QN(
        \xmem_inst/mem[19][31] ) );
  DFF_X1 \xmem_inst/mem_reg[19][30]  ( .D(n4782), .CK(clk), .QN(
        \xmem_inst/mem[19][30] ) );
  DFF_X1 \xmem_inst/mem_reg[19][19]  ( .D(n4771), .CK(clk), .QN(
        \xmem_inst/mem[19][19] ) );
  DFF_X1 \xmem_inst/mem_reg[19][15]  ( .D(n4767), .CK(clk), .QN(
        \xmem_inst/mem[19][15] ) );
  DFF_X1 \xmem_inst/mem_reg[18][31]  ( .D(n4751), .CK(clk), .QN(
        \xmem_inst/mem[18][31] ) );
  DFF_X1 \xmem_inst/mem_reg[18][30]  ( .D(n4750), .CK(clk), .QN(
        \xmem_inst/mem[18][30] ) );
  DFF_X1 \xmem_inst/mem_reg[18][19]  ( .D(n4739), .CK(clk), .QN(
        \xmem_inst/mem[18][19] ) );
  DFF_X1 \xmem_inst/mem_reg[18][15]  ( .D(n4735), .CK(clk), .QN(
        \xmem_inst/mem[18][15] ) );
  DFF_X1 \xmem_inst/mem_reg[17][31]  ( .D(n4719), .CK(clk), .QN(
        \xmem_inst/mem[17][31] ) );
  DFF_X1 \xmem_inst/mem_reg[17][30]  ( .D(n4718), .CK(clk), .QN(
        \xmem_inst/mem[17][30] ) );
  DFF_X1 \xmem_inst/mem_reg[17][19]  ( .D(n4707), .CK(clk), .QN(
        \xmem_inst/mem[17][19] ) );
  DFF_X1 \xmem_inst/mem_reg[17][15]  ( .D(n4703), .CK(clk), .QN(
        \xmem_inst/mem[17][15] ) );
  DFF_X1 \xmem_inst/mem_reg[16][31]  ( .D(n4687), .CK(clk), .QN(
        \xmem_inst/mem[16][31] ) );
  DFF_X1 \xmem_inst/mem_reg[16][30]  ( .D(n4686), .CK(clk), .QN(
        \xmem_inst/mem[16][30] ) );
  DFF_X1 \xmem_inst/mem_reg[16][19]  ( .D(n4675), .CK(clk), .QN(
        \xmem_inst/mem[16][19] ) );
  DFF_X1 \xmem_inst/mem_reg[16][15]  ( .D(n4671), .CK(clk), .QN(
        \xmem_inst/mem[16][15] ) );
  DFF_X1 \xmem_inst/mem_reg[7][31]  ( .D(n4399), .CK(clk), .QN(
        \xmem_inst/mem[7][31] ) );
  DFF_X1 \xmem_inst/mem_reg[7][30]  ( .D(n4398), .CK(clk), .QN(
        \xmem_inst/mem[7][30] ) );
  DFF_X1 \xmem_inst/mem_reg[7][19]  ( .D(n4388), .CK(clk), .QN(
        \xmem_inst/mem[7][19] ) );
  DFF_X1 \xmem_inst/mem_reg[7][15]  ( .D(n4384), .CK(clk), .QN(
        \xmem_inst/mem[7][15] ) );
  DFF_X1 \xmem_inst/mem_reg[6][31]  ( .D(n4368), .CK(clk), .QN(
        \xmem_inst/mem[6][31] ) );
  DFF_X1 \xmem_inst/mem_reg[6][30]  ( .D(n4367), .CK(clk), .QN(
        \xmem_inst/mem[6][30] ) );
  DFF_X1 \xmem_inst/mem_reg[6][19]  ( .D(n4356), .CK(clk), .QN(
        \xmem_inst/mem[6][19] ) );
  DFF_X1 \xmem_inst/mem_reg[6][15]  ( .D(n4352), .CK(clk), .QN(
        \xmem_inst/mem[6][15] ) );
  DFF_X1 \xmem_inst/mem_reg[5][31]  ( .D(n4336), .CK(clk), .QN(
        \xmem_inst/mem[5][31] ) );
  DFF_X1 \xmem_inst/mem_reg[5][30]  ( .D(n4335), .CK(clk), .QN(
        \xmem_inst/mem[5][30] ) );
  DFF_X1 \xmem_inst/mem_reg[5][19]  ( .D(n4324), .CK(clk), .QN(
        \xmem_inst/mem[5][19] ) );
  DFF_X1 \xmem_inst/mem_reg[5][15]  ( .D(n4320), .CK(clk), .QN(
        \xmem_inst/mem[5][15] ) );
  DFF_X1 \xmem_inst/mem_reg[4][31]  ( .D(n4304), .CK(clk), .QN(
        \xmem_inst/mem[4][31] ) );
  DFF_X1 \xmem_inst/mem_reg[4][30]  ( .D(n4303), .CK(clk), .QN(
        \xmem_inst/mem[4][30] ) );
  DFF_X1 \xmem_inst/mem_reg[4][19]  ( .D(n4292), .CK(clk), .QN(
        \xmem_inst/mem[4][19] ) );
  DFF_X1 \xmem_inst/mem_reg[4][15]  ( .D(n4288), .CK(clk), .QN(
        \xmem_inst/mem[4][15] ) );
  DFF_X1 \xmem_inst/mem_reg[3][31]  ( .D(n4272), .CK(clk), .QN(
        \xmem_inst/mem[3][31] ) );
  DFF_X1 \xmem_inst/mem_reg[3][30]  ( .D(n4271), .CK(clk), .QN(
        \xmem_inst/mem[3][30] ) );
  DFF_X1 \xmem_inst/mem_reg[3][19]  ( .D(n4260), .CK(clk), .QN(
        \xmem_inst/mem[3][19] ) );
  DFF_X1 \xmem_inst/mem_reg[3][15]  ( .D(n4256), .CK(clk), .QN(
        \xmem_inst/mem[3][15] ) );
  DFF_X1 \xmem_inst/mem_reg[2][31]  ( .D(n4240), .CK(clk), .QN(
        \xmem_inst/mem[2][31] ) );
  DFF_X1 \xmem_inst/mem_reg[2][30]  ( .D(n4239), .CK(clk), .QN(
        \xmem_inst/mem[2][30] ) );
  DFF_X1 \xmem_inst/mem_reg[2][19]  ( .D(n4228), .CK(clk), .QN(
        \xmem_inst/mem[2][19] ) );
  DFF_X1 \xmem_inst/mem_reg[2][15]  ( .D(n4224), .CK(clk), .QN(
        \xmem_inst/mem[2][15] ) );
  DFF_X1 \xmem_inst/mem_reg[1][31]  ( .D(n4208), .CK(clk), .QN(
        \xmem_inst/mem[1][31] ) );
  DFF_X1 \xmem_inst/mem_reg[1][30]  ( .D(n4207), .CK(clk), .QN(
        \xmem_inst/mem[1][30] ) );
  DFF_X1 \xmem_inst/mem_reg[1][19]  ( .D(n4196), .CK(clk), .QN(
        \xmem_inst/mem[1][19] ) );
  DFF_X1 \xmem_inst/mem_reg[1][15]  ( .D(n4192), .CK(clk), .QN(
        \xmem_inst/mem[1][15] ) );
  DFF_X1 \xmem_inst/mem_reg[0][31]  ( .D(n4176), .CK(clk), .QN(
        \xmem_inst/mem[0][31] ) );
  DFF_X1 \xmem_inst/mem_reg[0][30]  ( .D(n4175), .CK(clk), .QN(
        \xmem_inst/mem[0][30] ) );
  DFF_X1 \xmem_inst/mem_reg[0][19]  ( .D(n4164), .CK(clk), .QN(
        \xmem_inst/mem[0][19] ) );
  DFF_X1 \xmem_inst/mem_reg[0][15]  ( .D(n4160), .CK(clk), .QN(
        \xmem_inst/mem[0][15] ) );
  DFF_X1 \xmem_inst/mem_reg[23][29]  ( .D(n4909), .CK(clk), .QN(
        \xmem_inst/mem[23][29] ) );
  DFF_X1 \xmem_inst/mem_reg[23][27]  ( .D(n4907), .CK(clk), .QN(
        \xmem_inst/mem[23][27] ) );
  DFF_X1 \xmem_inst/mem_reg[23][25]  ( .D(n4905), .CK(clk), .QN(
        \xmem_inst/mem[23][25] ) );
  DFF_X1 \xmem_inst/mem_reg[23][14]  ( .D(n4894), .CK(clk), .QN(
        \xmem_inst/mem[23][14] ) );
  DFF_X1 \xmem_inst/mem_reg[23][11]  ( .D(n4891), .CK(clk), .QN(
        \xmem_inst/mem[23][11] ) );
  DFF_X1 \xmem_inst/mem_reg[23][9]  ( .D(n4889), .CK(clk), .QN(
        \xmem_inst/mem[23][9] ) );
  DFF_X1 \xmem_inst/mem_reg[23][8]  ( .D(n4888), .CK(clk), .QN(
        \xmem_inst/mem[23][8] ) );
  DFF_X1 \xmem_inst/mem_reg[23][7]  ( .D(n4887), .CK(clk), .QN(
        \xmem_inst/mem[23][7] ) );
  DFF_X1 \xmem_inst/mem_reg[23][6]  ( .D(n4886), .CK(clk), .QN(
        \xmem_inst/mem[23][6] ) );
  DFF_X1 \xmem_inst/mem_reg[23][5]  ( .D(n4885), .CK(clk), .QN(
        \xmem_inst/mem[23][5] ) );
  DFF_X1 \xmem_inst/mem_reg[22][29]  ( .D(n4877), .CK(clk), .QN(
        \xmem_inst/mem[22][29] ) );
  DFF_X1 \xmem_inst/mem_reg[22][27]  ( .D(n4875), .CK(clk), .QN(
        \xmem_inst/mem[22][27] ) );
  DFF_X1 \xmem_inst/mem_reg[22][25]  ( .D(n4873), .CK(clk), .QN(
        \xmem_inst/mem[22][25] ) );
  DFF_X1 \xmem_inst/mem_reg[22][14]  ( .D(n4862), .CK(clk), .QN(
        \xmem_inst/mem[22][14] ) );
  DFF_X1 \xmem_inst/mem_reg[22][11]  ( .D(n4859), .CK(clk), .QN(
        \xmem_inst/mem[22][11] ) );
  DFF_X1 \xmem_inst/mem_reg[22][9]  ( .D(n4857), .CK(clk), .QN(
        \xmem_inst/mem[22][9] ) );
  DFF_X1 \xmem_inst/mem_reg[22][8]  ( .D(n4856), .CK(clk), .QN(
        \xmem_inst/mem[22][8] ) );
  DFF_X1 \xmem_inst/mem_reg[22][7]  ( .D(n4855), .CK(clk), .QN(
        \xmem_inst/mem[22][7] ) );
  DFF_X1 \xmem_inst/mem_reg[22][6]  ( .D(n4854), .CK(clk), .QN(
        \xmem_inst/mem[22][6] ) );
  DFF_X1 \xmem_inst/mem_reg[22][5]  ( .D(n4853), .CK(clk), .QN(
        \xmem_inst/mem[22][5] ) );
  DFF_X1 \xmem_inst/mem_reg[21][29]  ( .D(n4845), .CK(clk), .QN(
        \xmem_inst/mem[21][29] ) );
  DFF_X1 \xmem_inst/mem_reg[21][27]  ( .D(n4843), .CK(clk), .QN(
        \xmem_inst/mem[21][27] ) );
  DFF_X1 \xmem_inst/mem_reg[21][25]  ( .D(n4841), .CK(clk), .QN(
        \xmem_inst/mem[21][25] ) );
  DFF_X1 \xmem_inst/mem_reg[21][14]  ( .D(n4830), .CK(clk), .QN(
        \xmem_inst/mem[21][14] ) );
  DFF_X1 \xmem_inst/mem_reg[21][11]  ( .D(n4827), .CK(clk), .QN(
        \xmem_inst/mem[21][11] ) );
  DFF_X1 \xmem_inst/mem_reg[21][9]  ( .D(n4825), .CK(clk), .QN(
        \xmem_inst/mem[21][9] ) );
  DFF_X1 \xmem_inst/mem_reg[21][8]  ( .D(n4824), .CK(clk), .QN(
        \xmem_inst/mem[21][8] ) );
  DFF_X1 \xmem_inst/mem_reg[21][7]  ( .D(n4823), .CK(clk), .QN(
        \xmem_inst/mem[21][7] ) );
  DFF_X1 \xmem_inst/mem_reg[21][6]  ( .D(n4822), .CK(clk), .QN(
        \xmem_inst/mem[21][6] ) );
  DFF_X1 \xmem_inst/mem_reg[21][5]  ( .D(n4821), .CK(clk), .QN(
        \xmem_inst/mem[21][5] ) );
  DFF_X1 \xmem_inst/mem_reg[20][29]  ( .D(n4813), .CK(clk), .QN(
        \xmem_inst/mem[20][29] ) );
  DFF_X1 \xmem_inst/mem_reg[20][27]  ( .D(n4811), .CK(clk), .QN(
        \xmem_inst/mem[20][27] ) );
  DFF_X1 \xmem_inst/mem_reg[20][25]  ( .D(n4809), .CK(clk), .QN(
        \xmem_inst/mem[20][25] ) );
  DFF_X1 \xmem_inst/mem_reg[20][14]  ( .D(n4798), .CK(clk), .QN(
        \xmem_inst/mem[20][14] ) );
  DFF_X1 \xmem_inst/mem_reg[20][11]  ( .D(n4795), .CK(clk), .QN(
        \xmem_inst/mem[20][11] ) );
  DFF_X1 \xmem_inst/mem_reg[20][9]  ( .D(n4793), .CK(clk), .QN(
        \xmem_inst/mem[20][9] ) );
  DFF_X1 \xmem_inst/mem_reg[20][8]  ( .D(n4792), .CK(clk), .QN(
        \xmem_inst/mem[20][8] ) );
  DFF_X1 \xmem_inst/mem_reg[20][7]  ( .D(n4791), .CK(clk), .QN(
        \xmem_inst/mem[20][7] ) );
  DFF_X1 \xmem_inst/mem_reg[20][6]  ( .D(n4790), .CK(clk), .QN(
        \xmem_inst/mem[20][6] ) );
  DFF_X1 \xmem_inst/mem_reg[20][5]  ( .D(n4789), .CK(clk), .QN(
        \xmem_inst/mem[20][5] ) );
  DFF_X1 \xmem_inst/mem_reg[7][29]  ( .D(n4397), .CK(clk), .QN(
        \xmem_inst/mem[7][29] ) );
  DFF_X1 \xmem_inst/mem_reg[7][27]  ( .D(n4395), .CK(clk), .QN(
        \xmem_inst/mem[7][27] ) );
  DFF_X1 \xmem_inst/mem_reg[7][25]  ( .D(n4393), .CK(clk), .QN(
        \xmem_inst/mem[7][25] ) );
  DFF_X1 \xmem_inst/mem_reg[7][14]  ( .D(n4383), .CK(clk), .QN(
        \xmem_inst/mem[7][14] ) );
  DFF_X1 \xmem_inst/mem_reg[7][11]  ( .D(n4380), .CK(clk), .QN(
        \xmem_inst/mem[7][11] ) );
  DFF_X1 \xmem_inst/mem_reg[7][9]  ( .D(n4378), .CK(clk), .QN(
        \xmem_inst/mem[7][9] ) );
  DFF_X1 \xmem_inst/mem_reg[7][7]  ( .D(n4376), .CK(clk), .QN(
        \xmem_inst/mem[7][7] ) );
  DFF_X1 \xmem_inst/mem_reg[7][6]  ( .D(n4375), .CK(clk), .QN(
        \xmem_inst/mem[7][6] ) );
  DFF_X1 \xmem_inst/mem_reg[7][5]  ( .D(n4374), .CK(clk), .QN(
        \xmem_inst/mem[7][5] ) );
  DFF_X1 \xmem_inst/mem_reg[6][29]  ( .D(n4366), .CK(clk), .QN(
        \xmem_inst/mem[6][29] ) );
  DFF_X1 \xmem_inst/mem_reg[6][27]  ( .D(n4364), .CK(clk), .QN(
        \xmem_inst/mem[6][27] ) );
  DFF_X1 \xmem_inst/mem_reg[6][25]  ( .D(n4362), .CK(clk), .QN(
        \xmem_inst/mem[6][25] ) );
  DFF_X1 \xmem_inst/mem_reg[6][14]  ( .D(n4351), .CK(clk), .QN(
        \xmem_inst/mem[6][14] ) );
  DFF_X1 \xmem_inst/mem_reg[6][11]  ( .D(n4348), .CK(clk), .QN(
        \xmem_inst/mem[6][11] ) );
  DFF_X1 \xmem_inst/mem_reg[6][9]  ( .D(n4346), .CK(clk), .QN(
        \xmem_inst/mem[6][9] ) );
  DFF_X1 \xmem_inst/mem_reg[6][8]  ( .D(n4345), .CK(clk), .QN(
        \xmem_inst/mem[6][8] ) );
  DFF_X1 \xmem_inst/mem_reg[6][7]  ( .D(n4344), .CK(clk), .QN(
        \xmem_inst/mem[6][7] ) );
  DFF_X1 \xmem_inst/mem_reg[6][6]  ( .D(n4343), .CK(clk), .QN(
        \xmem_inst/mem[6][6] ) );
  DFF_X1 \xmem_inst/mem_reg[6][5]  ( .D(n4342), .CK(clk), .QN(
        \xmem_inst/mem[6][5] ) );
  DFF_X1 \xmem_inst/mem_reg[5][29]  ( .D(n4334), .CK(clk), .QN(
        \xmem_inst/mem[5][29] ) );
  DFF_X1 \xmem_inst/mem_reg[5][27]  ( .D(n4332), .CK(clk), .QN(
        \xmem_inst/mem[5][27] ) );
  DFF_X1 \xmem_inst/mem_reg[5][25]  ( .D(n4330), .CK(clk), .QN(
        \xmem_inst/mem[5][25] ) );
  DFF_X1 \xmem_inst/mem_reg[5][14]  ( .D(n4319), .CK(clk), .QN(
        \xmem_inst/mem[5][14] ) );
  DFF_X1 \xmem_inst/mem_reg[5][11]  ( .D(n4316), .CK(clk), .QN(
        \xmem_inst/mem[5][11] ) );
  DFF_X1 \xmem_inst/mem_reg[5][9]  ( .D(n4314), .CK(clk), .QN(
        \xmem_inst/mem[5][9] ) );
  DFF_X1 \xmem_inst/mem_reg[5][8]  ( .D(n4313), .CK(clk), .QN(
        \xmem_inst/mem[5][8] ) );
  DFF_X1 \xmem_inst/mem_reg[5][7]  ( .D(n4312), .CK(clk), .QN(
        \xmem_inst/mem[5][7] ) );
  DFF_X1 \xmem_inst/mem_reg[5][6]  ( .D(n4311), .CK(clk), .QN(
        \xmem_inst/mem[5][6] ) );
  DFF_X1 \xmem_inst/mem_reg[5][5]  ( .D(n4310), .CK(clk), .QN(
        \xmem_inst/mem[5][5] ) );
  DFF_X1 \xmem_inst/mem_reg[4][29]  ( .D(n4302), .CK(clk), .QN(
        \xmem_inst/mem[4][29] ) );
  DFF_X1 \xmem_inst/mem_reg[4][27]  ( .D(n4300), .CK(clk), .QN(
        \xmem_inst/mem[4][27] ) );
  DFF_X1 \xmem_inst/mem_reg[4][25]  ( .D(n4298), .CK(clk), .QN(
        \xmem_inst/mem[4][25] ) );
  DFF_X1 \xmem_inst/mem_reg[4][14]  ( .D(n4287), .CK(clk), .QN(
        \xmem_inst/mem[4][14] ) );
  DFF_X1 \xmem_inst/mem_reg[4][11]  ( .D(n4284), .CK(clk), .QN(
        \xmem_inst/mem[4][11] ) );
  DFF_X1 \xmem_inst/mem_reg[4][9]  ( .D(n4282), .CK(clk), .QN(
        \xmem_inst/mem[4][9] ) );
  DFF_X1 \xmem_inst/mem_reg[4][8]  ( .D(n4281), .CK(clk), .QN(
        \xmem_inst/mem[4][8] ) );
  DFF_X1 \xmem_inst/mem_reg[4][7]  ( .D(n4280), .CK(clk), .QN(
        \xmem_inst/mem[4][7] ) );
  DFF_X1 \xmem_inst/mem_reg[4][6]  ( .D(n4279), .CK(clk), .QN(
        \xmem_inst/mem[4][6] ) );
  DFF_X1 \xmem_inst/mem_reg[4][5]  ( .D(n4278), .CK(clk), .QN(
        \xmem_inst/mem[4][5] ) );
  DFF_X1 \xmem_inst/mem_reg[19][29]  ( .D(n4781), .CK(clk), .QN(
        \xmem_inst/mem[19][29] ) );
  DFF_X1 \xmem_inst/mem_reg[19][27]  ( .D(n4779), .CK(clk), .QN(
        \xmem_inst/mem[19][27] ) );
  DFF_X1 \xmem_inst/mem_reg[19][25]  ( .D(n4777), .CK(clk), .QN(
        \xmem_inst/mem[19][25] ) );
  DFF_X1 \xmem_inst/mem_reg[19][14]  ( .D(n4766), .CK(clk), .QN(
        \xmem_inst/mem[19][14] ) );
  DFF_X1 \xmem_inst/mem_reg[19][11]  ( .D(n4763), .CK(clk), .QN(
        \xmem_inst/mem[19][11] ) );
  DFF_X1 \xmem_inst/mem_reg[19][9]  ( .D(n4761), .CK(clk), .QN(
        \xmem_inst/mem[19][9] ) );
  DFF_X1 \xmem_inst/mem_reg[19][8]  ( .D(n4760), .CK(clk), .QN(
        \xmem_inst/mem[19][8] ) );
  DFF_X1 \xmem_inst/mem_reg[19][7]  ( .D(n4759), .CK(clk), .QN(
        \xmem_inst/mem[19][7] ) );
  DFF_X1 \xmem_inst/mem_reg[19][6]  ( .D(n4758), .CK(clk), .QN(
        \xmem_inst/mem[19][6] ) );
  DFF_X1 \xmem_inst/mem_reg[19][5]  ( .D(n4757), .CK(clk), .QN(
        \xmem_inst/mem[19][5] ) );
  DFF_X1 \xmem_inst/mem_reg[3][29]  ( .D(n4270), .CK(clk), .QN(
        \xmem_inst/mem[3][29] ) );
  DFF_X1 \xmem_inst/mem_reg[3][27]  ( .D(n4268), .CK(clk), .QN(
        \xmem_inst/mem[3][27] ) );
  DFF_X1 \xmem_inst/mem_reg[3][25]  ( .D(n4266), .CK(clk), .QN(
        \xmem_inst/mem[3][25] ) );
  DFF_X1 \xmem_inst/mem_reg[3][14]  ( .D(n4255), .CK(clk), .QN(
        \xmem_inst/mem[3][14] ) );
  DFF_X1 \xmem_inst/mem_reg[3][11]  ( .D(n4252), .CK(clk), .QN(
        \xmem_inst/mem[3][11] ) );
  DFF_X1 \xmem_inst/mem_reg[3][9]  ( .D(n4250), .CK(clk), .QN(
        \xmem_inst/mem[3][9] ) );
  DFF_X1 \xmem_inst/mem_reg[3][8]  ( .D(n4249), .CK(clk), .QN(
        \xmem_inst/mem[3][8] ) );
  DFF_X1 \xmem_inst/mem_reg[3][7]  ( .D(n4248), .CK(clk), .QN(
        \xmem_inst/mem[3][7] ) );
  DFF_X1 \xmem_inst/mem_reg[3][6]  ( .D(n4247), .CK(clk), .QN(
        \xmem_inst/mem[3][6] ) );
  DFF_X1 \xmem_inst/mem_reg[3][5]  ( .D(n4246), .CK(clk), .QN(
        \xmem_inst/mem[3][5] ) );
  DFF_X1 \xmem_inst/mem_reg[23][28]  ( .D(n4908), .CK(clk), .QN(
        \xmem_inst/mem[23][28] ) );
  DFF_X1 \xmem_inst/mem_reg[23][26]  ( .D(n4906), .CK(clk), .QN(
        \xmem_inst/mem[23][26] ) );
  DFF_X1 \xmem_inst/mem_reg[23][24]  ( .D(n4904), .CK(clk), .QN(
        \xmem_inst/mem[23][24] ) );
  DFF_X1 \xmem_inst/mem_reg[23][23]  ( .D(n4903), .CK(clk), .QN(
        \xmem_inst/mem[23][23] ) );
  DFF_X1 \xmem_inst/mem_reg[23][22]  ( .D(n4902), .CK(clk), .QN(
        \xmem_inst/mem[23][22] ) );
  DFF_X1 \xmem_inst/mem_reg[23][21]  ( .D(n4901), .CK(clk), .QN(
        \xmem_inst/mem[23][21] ) );
  DFF_X1 \xmem_inst/mem_reg[23][20]  ( .D(n4900), .CK(clk), .QN(
        \xmem_inst/mem[23][20] ) );
  DFF_X1 \xmem_inst/mem_reg[23][18]  ( .D(n4898), .CK(clk), .QN(
        \xmem_inst/mem[23][18] ) );
  DFF_X1 \xmem_inst/mem_reg[23][17]  ( .D(n4897), .CK(clk), .QN(
        \xmem_inst/mem[23][17] ) );
  DFF_X1 \xmem_inst/mem_reg[23][16]  ( .D(n4896), .CK(clk), .QN(
        \xmem_inst/mem[23][16] ) );
  DFF_X1 \xmem_inst/mem_reg[23][13]  ( .D(n4893), .CK(clk), .QN(
        \xmem_inst/mem[23][13] ) );
  DFF_X1 \xmem_inst/mem_reg[23][12]  ( .D(n4892), .CK(clk), .QN(
        \xmem_inst/mem[23][12] ) );
  DFF_X1 \xmem_inst/mem_reg[23][10]  ( .D(n4890), .CK(clk), .QN(
        \xmem_inst/mem[23][10] ) );
  DFF_X1 \xmem_inst/mem_reg[23][4]  ( .D(n4884), .CK(clk), .QN(
        \xmem_inst/mem[23][4] ) );
  DFF_X1 \xmem_inst/mem_reg[23][3]  ( .D(n4883), .CK(clk), .QN(
        \xmem_inst/mem[23][3] ) );
  DFF_X1 \xmem_inst/mem_reg[23][2]  ( .D(n4882), .CK(clk), .QN(
        \xmem_inst/mem[23][2] ) );
  DFF_X1 \xmem_inst/mem_reg[23][1]  ( .D(n4881), .CK(clk), .QN(
        \xmem_inst/mem[23][1] ) );
  DFF_X1 \xmem_inst/mem_reg[23][0]  ( .D(n4880), .CK(clk), .QN(
        \xmem_inst/mem[23][0] ) );
  DFF_X1 \xmem_inst/mem_reg[22][28]  ( .D(n4876), .CK(clk), .QN(
        \xmem_inst/mem[22][28] ) );
  DFF_X1 \xmem_inst/mem_reg[22][26]  ( .D(n4874), .CK(clk), .QN(
        \xmem_inst/mem[22][26] ) );
  DFF_X1 \xmem_inst/mem_reg[22][24]  ( .D(n4872), .CK(clk), .QN(
        \xmem_inst/mem[22][24] ) );
  DFF_X1 \xmem_inst/mem_reg[22][23]  ( .D(n4871), .CK(clk), .QN(
        \xmem_inst/mem[22][23] ) );
  DFF_X1 \xmem_inst/mem_reg[22][22]  ( .D(n4870), .CK(clk), .QN(
        \xmem_inst/mem[22][22] ) );
  DFF_X1 \xmem_inst/mem_reg[22][21]  ( .D(n4869), .CK(clk), .QN(
        \xmem_inst/mem[22][21] ) );
  DFF_X1 \xmem_inst/mem_reg[22][20]  ( .D(n4868), .CK(clk), .QN(
        \xmem_inst/mem[22][20] ) );
  DFF_X1 \xmem_inst/mem_reg[22][18]  ( .D(n4866), .CK(clk), .QN(
        \xmem_inst/mem[22][18] ) );
  DFF_X1 \xmem_inst/mem_reg[22][17]  ( .D(n4865), .CK(clk), .QN(
        \xmem_inst/mem[22][17] ) );
  DFF_X1 \xmem_inst/mem_reg[22][16]  ( .D(n4864), .CK(clk), .QN(
        \xmem_inst/mem[22][16] ) );
  DFF_X1 \xmem_inst/mem_reg[22][13]  ( .D(n4861), .CK(clk), .QN(
        \xmem_inst/mem[22][13] ) );
  DFF_X1 \xmem_inst/mem_reg[22][12]  ( .D(n4860), .CK(clk), .QN(
        \xmem_inst/mem[22][12] ) );
  DFF_X1 \xmem_inst/mem_reg[22][10]  ( .D(n4858), .CK(clk), .QN(
        \xmem_inst/mem[22][10] ) );
  DFF_X1 \xmem_inst/mem_reg[22][4]  ( .D(n4852), .CK(clk), .QN(
        \xmem_inst/mem[22][4] ) );
  DFF_X1 \xmem_inst/mem_reg[22][3]  ( .D(n4851), .CK(clk), .QN(
        \xmem_inst/mem[22][3] ) );
  DFF_X1 \xmem_inst/mem_reg[22][2]  ( .D(n4850), .CK(clk), .QN(
        \xmem_inst/mem[22][2] ) );
  DFF_X1 \xmem_inst/mem_reg[22][1]  ( .D(n4849), .CK(clk), .QN(
        \xmem_inst/mem[22][1] ) );
  DFF_X1 \xmem_inst/mem_reg[22][0]  ( .D(n4848), .CK(clk), .QN(
        \xmem_inst/mem[22][0] ) );
  DFF_X1 \xmem_inst/mem_reg[21][28]  ( .D(n4844), .CK(clk), .QN(
        \xmem_inst/mem[21][28] ) );
  DFF_X1 \xmem_inst/mem_reg[21][26]  ( .D(n4842), .CK(clk), .QN(
        \xmem_inst/mem[21][26] ) );
  DFF_X1 \xmem_inst/mem_reg[21][24]  ( .D(n4840), .CK(clk), .QN(
        \xmem_inst/mem[21][24] ) );
  DFF_X1 \xmem_inst/mem_reg[21][23]  ( .D(n4839), .CK(clk), .QN(
        \xmem_inst/mem[21][23] ) );
  DFF_X1 \xmem_inst/mem_reg[21][22]  ( .D(n4838), .CK(clk), .QN(
        \xmem_inst/mem[21][22] ) );
  DFF_X1 \xmem_inst/mem_reg[21][21]  ( .D(n4837), .CK(clk), .QN(
        \xmem_inst/mem[21][21] ) );
  DFF_X1 \xmem_inst/mem_reg[21][20]  ( .D(n4836), .CK(clk), .QN(
        \xmem_inst/mem[21][20] ) );
  DFF_X1 \xmem_inst/mem_reg[21][18]  ( .D(n4834), .CK(clk), .QN(
        \xmem_inst/mem[21][18] ) );
  DFF_X1 \xmem_inst/mem_reg[21][17]  ( .D(n4833), .CK(clk), .QN(
        \xmem_inst/mem[21][17] ) );
  DFF_X1 \xmem_inst/mem_reg[21][16]  ( .D(n4832), .CK(clk), .QN(
        \xmem_inst/mem[21][16] ) );
  DFF_X1 \xmem_inst/mem_reg[21][13]  ( .D(n4829), .CK(clk), .QN(
        \xmem_inst/mem[21][13] ) );
  DFF_X1 \xmem_inst/mem_reg[21][12]  ( .D(n4828), .CK(clk), .QN(
        \xmem_inst/mem[21][12] ) );
  DFF_X1 \xmem_inst/mem_reg[21][10]  ( .D(n4826), .CK(clk), .QN(
        \xmem_inst/mem[21][10] ) );
  DFF_X1 \xmem_inst/mem_reg[21][4]  ( .D(n4820), .CK(clk), .QN(
        \xmem_inst/mem[21][4] ) );
  DFF_X1 \xmem_inst/mem_reg[21][3]  ( .D(n4819), .CK(clk), .QN(
        \xmem_inst/mem[21][3] ) );
  DFF_X1 \xmem_inst/mem_reg[21][2]  ( .D(n4818), .CK(clk), .QN(
        \xmem_inst/mem[21][2] ) );
  DFF_X1 \xmem_inst/mem_reg[21][1]  ( .D(n4817), .CK(clk), .QN(
        \xmem_inst/mem[21][1] ) );
  DFF_X1 \xmem_inst/mem_reg[21][0]  ( .D(n4816), .CK(clk), .QN(
        \xmem_inst/mem[21][0] ) );
  DFF_X1 \xmem_inst/mem_reg[20][28]  ( .D(n4812), .CK(clk), .QN(
        \xmem_inst/mem[20][28] ) );
  DFF_X1 \xmem_inst/mem_reg[20][26]  ( .D(n4810), .CK(clk), .QN(
        \xmem_inst/mem[20][26] ) );
  DFF_X1 \xmem_inst/mem_reg[20][24]  ( .D(n4808), .CK(clk), .QN(
        \xmem_inst/mem[20][24] ) );
  DFF_X1 \xmem_inst/mem_reg[20][23]  ( .D(n4807), .CK(clk), .QN(
        \xmem_inst/mem[20][23] ) );
  DFF_X1 \xmem_inst/mem_reg[20][22]  ( .D(n4806), .CK(clk), .QN(
        \xmem_inst/mem[20][22] ) );
  DFF_X1 \xmem_inst/mem_reg[20][21]  ( .D(n4805), .CK(clk), .QN(
        \xmem_inst/mem[20][21] ) );
  DFF_X1 \xmem_inst/mem_reg[20][20]  ( .D(n4804), .CK(clk), .QN(
        \xmem_inst/mem[20][20] ) );
  DFF_X1 \xmem_inst/mem_reg[20][18]  ( .D(n4802), .CK(clk), .QN(
        \xmem_inst/mem[20][18] ) );
  DFF_X1 \xmem_inst/mem_reg[20][17]  ( .D(n4801), .CK(clk), .QN(
        \xmem_inst/mem[20][17] ) );
  DFF_X1 \xmem_inst/mem_reg[20][16]  ( .D(n4800), .CK(clk), .QN(
        \xmem_inst/mem[20][16] ) );
  DFF_X1 \xmem_inst/mem_reg[20][13]  ( .D(n4797), .CK(clk), .QN(
        \xmem_inst/mem[20][13] ) );
  DFF_X1 \xmem_inst/mem_reg[20][12]  ( .D(n4796), .CK(clk), .QN(
        \xmem_inst/mem[20][12] ) );
  DFF_X1 \xmem_inst/mem_reg[20][10]  ( .D(n4794), .CK(clk), .QN(
        \xmem_inst/mem[20][10] ) );
  DFF_X1 \xmem_inst/mem_reg[20][4]  ( .D(n4788), .CK(clk), .QN(
        \xmem_inst/mem[20][4] ) );
  DFF_X1 \xmem_inst/mem_reg[20][3]  ( .D(n4787), .CK(clk), .QN(
        \xmem_inst/mem[20][3] ) );
  DFF_X1 \xmem_inst/mem_reg[20][2]  ( .D(n4786), .CK(clk), .QN(
        \xmem_inst/mem[20][2] ) );
  DFF_X1 \xmem_inst/mem_reg[20][1]  ( .D(n4785), .CK(clk), .QN(
        \xmem_inst/mem[20][1] ) );
  DFF_X1 \xmem_inst/mem_reg[20][0]  ( .D(n4784), .CK(clk), .QN(
        \xmem_inst/mem[20][0] ) );
  DFF_X1 \xmem_inst/mem_reg[19][28]  ( .D(n4780), .CK(clk), .QN(
        \xmem_inst/mem[19][28] ) );
  DFF_X1 \xmem_inst/mem_reg[19][26]  ( .D(n4778), .CK(clk), .QN(
        \xmem_inst/mem[19][26] ) );
  DFF_X1 \xmem_inst/mem_reg[19][24]  ( .D(n4776), .CK(clk), .QN(
        \xmem_inst/mem[19][24] ) );
  DFF_X1 \xmem_inst/mem_reg[19][23]  ( .D(n4775), .CK(clk), .QN(
        \xmem_inst/mem[19][23] ) );
  DFF_X1 \xmem_inst/mem_reg[19][22]  ( .D(n4774), .CK(clk), .QN(
        \xmem_inst/mem[19][22] ) );
  DFF_X1 \xmem_inst/mem_reg[19][21]  ( .D(n4773), .CK(clk), .QN(
        \xmem_inst/mem[19][21] ) );
  DFF_X1 \xmem_inst/mem_reg[19][20]  ( .D(n4772), .CK(clk), .QN(
        \xmem_inst/mem[19][20] ) );
  DFF_X1 \xmem_inst/mem_reg[19][18]  ( .D(n4770), .CK(clk), .QN(
        \xmem_inst/mem[19][18] ) );
  DFF_X1 \xmem_inst/mem_reg[19][17]  ( .D(n4769), .CK(clk), .QN(
        \xmem_inst/mem[19][17] ) );
  DFF_X1 \xmem_inst/mem_reg[19][16]  ( .D(n4768), .CK(clk), .QN(
        \xmem_inst/mem[19][16] ) );
  DFF_X1 \xmem_inst/mem_reg[19][13]  ( .D(n4765), .CK(clk), .QN(
        \xmem_inst/mem[19][13] ) );
  DFF_X1 \xmem_inst/mem_reg[19][12]  ( .D(n4764), .CK(clk), .QN(
        \xmem_inst/mem[19][12] ) );
  DFF_X1 \xmem_inst/mem_reg[19][10]  ( .D(n4762), .CK(clk), .QN(
        \xmem_inst/mem[19][10] ) );
  DFF_X1 \xmem_inst/mem_reg[19][4]  ( .D(n4756), .CK(clk), .QN(
        \xmem_inst/mem[19][4] ) );
  DFF_X1 \xmem_inst/mem_reg[19][3]  ( .D(n4755), .CK(clk), .QN(
        \xmem_inst/mem[19][3] ) );
  DFF_X1 \xmem_inst/mem_reg[19][2]  ( .D(n4754), .CK(clk), .QN(
        \xmem_inst/mem[19][2] ) );
  DFF_X1 \xmem_inst/mem_reg[19][1]  ( .D(n4753), .CK(clk), .QN(
        \xmem_inst/mem[19][1] ) );
  DFF_X1 \xmem_inst/mem_reg[19][0]  ( .D(n4752), .CK(clk), .QN(
        \xmem_inst/mem[19][0] ) );
  DFF_X1 \xmem_inst/mem_reg[18][28]  ( .D(n4748), .CK(clk), .QN(
        \xmem_inst/mem[18][28] ) );
  DFF_X1 \xmem_inst/mem_reg[18][26]  ( .D(n4746), .CK(clk), .QN(
        \xmem_inst/mem[18][26] ) );
  DFF_X1 \xmem_inst/mem_reg[18][24]  ( .D(n4744), .CK(clk), .QN(
        \xmem_inst/mem[18][24] ) );
  DFF_X1 \xmem_inst/mem_reg[18][23]  ( .D(n4743), .CK(clk), .QN(
        \xmem_inst/mem[18][23] ) );
  DFF_X1 \xmem_inst/mem_reg[18][22]  ( .D(n4742), .CK(clk), .QN(
        \xmem_inst/mem[18][22] ) );
  DFF_X1 \xmem_inst/mem_reg[18][21]  ( .D(n4741), .CK(clk), .QN(
        \xmem_inst/mem[18][21] ) );
  DFF_X1 \xmem_inst/mem_reg[18][20]  ( .D(n4740), .CK(clk), .QN(
        \xmem_inst/mem[18][20] ) );
  DFF_X1 \xmem_inst/mem_reg[18][18]  ( .D(n4738), .CK(clk), .QN(
        \xmem_inst/mem[18][18] ) );
  DFF_X1 \xmem_inst/mem_reg[18][17]  ( .D(n4737), .CK(clk), .QN(
        \xmem_inst/mem[18][17] ) );
  DFF_X1 \xmem_inst/mem_reg[18][16]  ( .D(n4736), .CK(clk), .QN(
        \xmem_inst/mem[18][16] ) );
  DFF_X1 \xmem_inst/mem_reg[18][13]  ( .D(n4733), .CK(clk), .QN(
        \xmem_inst/mem[18][13] ) );
  DFF_X1 \xmem_inst/mem_reg[18][12]  ( .D(n4732), .CK(clk), .QN(
        \xmem_inst/mem[18][12] ) );
  DFF_X1 \xmem_inst/mem_reg[18][10]  ( .D(n4730), .CK(clk), .QN(
        \xmem_inst/mem[18][10] ) );
  DFF_X1 \xmem_inst/mem_reg[18][4]  ( .D(n4724), .CK(clk), .QN(
        \xmem_inst/mem[18][4] ) );
  DFF_X1 \xmem_inst/mem_reg[18][3]  ( .D(n4723), .CK(clk), .QN(
        \xmem_inst/mem[18][3] ) );
  DFF_X1 \xmem_inst/mem_reg[18][2]  ( .D(n4722), .CK(clk), .QN(
        \xmem_inst/mem[18][2] ) );
  DFF_X1 \xmem_inst/mem_reg[18][1]  ( .D(n4721), .CK(clk), .QN(
        \xmem_inst/mem[18][1] ) );
  DFF_X1 \xmem_inst/mem_reg[18][0]  ( .D(n4720), .CK(clk), .QN(
        \xmem_inst/mem[18][0] ) );
  DFF_X1 \xmem_inst/mem_reg[7][28]  ( .D(n4396), .CK(clk), .QN(
        \xmem_inst/mem[7][28] ) );
  DFF_X1 \xmem_inst/mem_reg[7][26]  ( .D(n4394), .CK(clk), .QN(
        \xmem_inst/mem[7][26] ) );
  DFF_X1 \xmem_inst/mem_reg[7][24]  ( .D(n4392), .CK(clk), .QN(
        \xmem_inst/mem[7][24] ) );
  DFF_X1 \xmem_inst/mem_reg[7][23]  ( .D(n4391), .CK(clk), .QN(
        \xmem_inst/mem[7][23] ) );
  DFF_X1 \xmem_inst/mem_reg[7][22]  ( .D(n4390), .CK(clk), .QN(
        \xmem_inst/mem[7][22] ) );
  DFF_X1 \xmem_inst/mem_reg[7][21]  ( .D(n4389), .CK(clk), .QN(
        \xmem_inst/mem[7][21] ) );
  DFF_X1 \xmem_inst/mem_reg[7][18]  ( .D(n4387), .CK(clk), .QN(
        \xmem_inst/mem[7][18] ) );
  DFF_X1 \xmem_inst/mem_reg[7][17]  ( .D(n4386), .CK(clk), .QN(
        \xmem_inst/mem[7][17] ) );
  DFF_X1 \xmem_inst/mem_reg[7][16]  ( .D(n4385), .CK(clk), .QN(
        \xmem_inst/mem[7][16] ) );
  DFF_X1 \xmem_inst/mem_reg[7][13]  ( .D(n4382), .CK(clk), .QN(
        \xmem_inst/mem[7][13] ) );
  DFF_X1 \xmem_inst/mem_reg[7][12]  ( .D(n4381), .CK(clk), .QN(
        \xmem_inst/mem[7][12] ) );
  DFF_X1 \xmem_inst/mem_reg[7][10]  ( .D(n4379), .CK(clk), .QN(
        \xmem_inst/mem[7][10] ) );
  DFF_X1 \xmem_inst/mem_reg[7][4]  ( .D(n4373), .CK(clk), .QN(
        \xmem_inst/mem[7][4] ) );
  DFF_X1 \xmem_inst/mem_reg[7][3]  ( .D(n4372), .CK(clk), .QN(
        \xmem_inst/mem[7][3] ) );
  DFF_X1 \xmem_inst/mem_reg[7][2]  ( .D(n4371), .CK(clk), .QN(
        \xmem_inst/mem[7][2] ) );
  DFF_X1 \xmem_inst/mem_reg[7][1]  ( .D(n4370), .CK(clk), .QN(
        \xmem_inst/mem[7][1] ) );
  DFF_X1 \xmem_inst/mem_reg[7][0]  ( .D(n4369), .CK(clk), .QN(
        \xmem_inst/mem[7][0] ) );
  DFF_X1 \xmem_inst/mem_reg[6][28]  ( .D(n4365), .CK(clk), .QN(
        \xmem_inst/mem[6][28] ) );
  DFF_X1 \xmem_inst/mem_reg[6][26]  ( .D(n4363), .CK(clk), .QN(
        \xmem_inst/mem[6][26] ) );
  DFF_X1 \xmem_inst/mem_reg[6][24]  ( .D(n4361), .CK(clk), .QN(
        \xmem_inst/mem[6][24] ) );
  DFF_X1 \xmem_inst/mem_reg[6][23]  ( .D(n4360), .CK(clk), .QN(
        \xmem_inst/mem[6][23] ) );
  DFF_X1 \xmem_inst/mem_reg[6][22]  ( .D(n4359), .CK(clk), .QN(
        \xmem_inst/mem[6][22] ) );
  DFF_X1 \xmem_inst/mem_reg[6][21]  ( .D(n4358), .CK(clk), .QN(
        \xmem_inst/mem[6][21] ) );
  DFF_X1 \xmem_inst/mem_reg[6][20]  ( .D(n4357), .CK(clk), .QN(
        \xmem_inst/mem[6][20] ) );
  DFF_X1 \xmem_inst/mem_reg[6][18]  ( .D(n4355), .CK(clk), .QN(
        \xmem_inst/mem[6][18] ) );
  DFF_X1 \xmem_inst/mem_reg[6][17]  ( .D(n4354), .CK(clk), .QN(
        \xmem_inst/mem[6][17] ) );
  DFF_X1 \xmem_inst/mem_reg[6][16]  ( .D(n4353), .CK(clk), .QN(
        \xmem_inst/mem[6][16] ) );
  DFF_X1 \xmem_inst/mem_reg[6][13]  ( .D(n4350), .CK(clk), .QN(
        \xmem_inst/mem[6][13] ) );
  DFF_X1 \xmem_inst/mem_reg[6][12]  ( .D(n4349), .CK(clk), .QN(
        \xmem_inst/mem[6][12] ) );
  DFF_X1 \xmem_inst/mem_reg[6][10]  ( .D(n4347), .CK(clk), .QN(
        \xmem_inst/mem[6][10] ) );
  DFF_X1 \xmem_inst/mem_reg[6][4]  ( .D(n4341), .CK(clk), .QN(
        \xmem_inst/mem[6][4] ) );
  DFF_X1 \xmem_inst/mem_reg[6][3]  ( .D(n4340), .CK(clk), .QN(
        \xmem_inst/mem[6][3] ) );
  DFF_X1 \xmem_inst/mem_reg[6][2]  ( .D(n4339), .CK(clk), .QN(
        \xmem_inst/mem[6][2] ) );
  DFF_X1 \xmem_inst/mem_reg[6][1]  ( .D(n4338), .CK(clk), .QN(
        \xmem_inst/mem[6][1] ) );
  DFF_X1 \xmem_inst/mem_reg[6][0]  ( .D(n4337), .CK(clk), .QN(
        \xmem_inst/mem[6][0] ) );
  DFF_X1 \xmem_inst/mem_reg[5][28]  ( .D(n4333), .CK(clk), .QN(
        \xmem_inst/mem[5][28] ) );
  DFF_X1 \xmem_inst/mem_reg[5][26]  ( .D(n4331), .CK(clk), .QN(
        \xmem_inst/mem[5][26] ) );
  DFF_X1 \xmem_inst/mem_reg[5][24]  ( .D(n4329), .CK(clk), .QN(
        \xmem_inst/mem[5][24] ) );
  DFF_X1 \xmem_inst/mem_reg[5][23]  ( .D(n4328), .CK(clk), .QN(
        \xmem_inst/mem[5][23] ) );
  DFF_X1 \xmem_inst/mem_reg[5][22]  ( .D(n4327), .CK(clk), .QN(
        \xmem_inst/mem[5][22] ) );
  DFF_X1 \xmem_inst/mem_reg[5][21]  ( .D(n4326), .CK(clk), .QN(
        \xmem_inst/mem[5][21] ) );
  DFF_X1 \xmem_inst/mem_reg[5][20]  ( .D(n4325), .CK(clk), .QN(
        \xmem_inst/mem[5][20] ) );
  DFF_X1 \xmem_inst/mem_reg[5][18]  ( .D(n4323), .CK(clk), .QN(
        \xmem_inst/mem[5][18] ) );
  DFF_X1 \xmem_inst/mem_reg[5][17]  ( .D(n4322), .CK(clk), .QN(
        \xmem_inst/mem[5][17] ) );
  DFF_X1 \xmem_inst/mem_reg[5][16]  ( .D(n4321), .CK(clk), .QN(
        \xmem_inst/mem[5][16] ) );
  DFF_X1 \xmem_inst/mem_reg[5][13]  ( .D(n4318), .CK(clk), .QN(
        \xmem_inst/mem[5][13] ) );
  DFF_X1 \xmem_inst/mem_reg[5][12]  ( .D(n4317), .CK(clk), .QN(
        \xmem_inst/mem[5][12] ) );
  DFF_X1 \xmem_inst/mem_reg[5][10]  ( .D(n4315), .CK(clk), .QN(
        \xmem_inst/mem[5][10] ) );
  DFF_X1 \xmem_inst/mem_reg[5][4]  ( .D(n4309), .CK(clk), .QN(
        \xmem_inst/mem[5][4] ) );
  DFF_X1 \xmem_inst/mem_reg[5][3]  ( .D(n4308), .CK(clk), .QN(
        \xmem_inst/mem[5][3] ) );
  DFF_X1 \xmem_inst/mem_reg[5][2]  ( .D(n4307), .CK(clk), .QN(
        \xmem_inst/mem[5][2] ) );
  DFF_X1 \xmem_inst/mem_reg[5][1]  ( .D(n4306), .CK(clk), .QN(
        \xmem_inst/mem[5][1] ) );
  DFF_X1 \xmem_inst/mem_reg[5][0]  ( .D(n4305), .CK(clk), .QN(
        \xmem_inst/mem[5][0] ) );
  DFF_X1 \xmem_inst/mem_reg[4][28]  ( .D(n4301), .CK(clk), .QN(
        \xmem_inst/mem[4][28] ) );
  DFF_X1 \xmem_inst/mem_reg[4][26]  ( .D(n4299), .CK(clk), .QN(
        \xmem_inst/mem[4][26] ) );
  DFF_X1 \xmem_inst/mem_reg[4][24]  ( .D(n4297), .CK(clk), .QN(
        \xmem_inst/mem[4][24] ) );
  DFF_X1 \xmem_inst/mem_reg[4][23]  ( .D(n4296), .CK(clk), .QN(
        \xmem_inst/mem[4][23] ) );
  DFF_X1 \xmem_inst/mem_reg[4][22]  ( .D(n4295), .CK(clk), .QN(
        \xmem_inst/mem[4][22] ) );
  DFF_X1 \xmem_inst/mem_reg[4][21]  ( .D(n4294), .CK(clk), .QN(
        \xmem_inst/mem[4][21] ) );
  DFF_X1 \xmem_inst/mem_reg[4][20]  ( .D(n4293), .CK(clk), .QN(
        \xmem_inst/mem[4][20] ) );
  DFF_X1 \xmem_inst/mem_reg[4][18]  ( .D(n4291), .CK(clk), .QN(
        \xmem_inst/mem[4][18] ) );
  DFF_X1 \xmem_inst/mem_reg[4][17]  ( .D(n4290), .CK(clk), .QN(
        \xmem_inst/mem[4][17] ) );
  DFF_X1 \xmem_inst/mem_reg[4][16]  ( .D(n4289), .CK(clk), .QN(
        \xmem_inst/mem[4][16] ) );
  DFF_X1 \xmem_inst/mem_reg[4][13]  ( .D(n4286), .CK(clk), .QN(
        \xmem_inst/mem[4][13] ) );
  DFF_X1 \xmem_inst/mem_reg[4][12]  ( .D(n4285), .CK(clk), .QN(
        \xmem_inst/mem[4][12] ) );
  DFF_X1 \xmem_inst/mem_reg[4][10]  ( .D(n4283), .CK(clk), .QN(
        \xmem_inst/mem[4][10] ) );
  DFF_X1 \xmem_inst/mem_reg[4][4]  ( .D(n4277), .CK(clk), .QN(
        \xmem_inst/mem[4][4] ) );
  DFF_X1 \xmem_inst/mem_reg[4][3]  ( .D(n4276), .CK(clk), .QN(
        \xmem_inst/mem[4][3] ) );
  DFF_X1 \xmem_inst/mem_reg[4][2]  ( .D(n4275), .CK(clk), .QN(
        \xmem_inst/mem[4][2] ) );
  DFF_X1 \xmem_inst/mem_reg[4][1]  ( .D(n4274), .CK(clk), .QN(
        \xmem_inst/mem[4][1] ) );
  DFF_X1 \xmem_inst/mem_reg[4][0]  ( .D(n4273), .CK(clk), .QN(
        \xmem_inst/mem[4][0] ) );
  DFF_X1 \xmem_inst/mem_reg[3][28]  ( .D(n4269), .CK(clk), .QN(
        \xmem_inst/mem[3][28] ) );
  DFF_X1 \xmem_inst/mem_reg[3][26]  ( .D(n4267), .CK(clk), .QN(
        \xmem_inst/mem[3][26] ) );
  DFF_X1 \xmem_inst/mem_reg[3][24]  ( .D(n4265), .CK(clk), .QN(
        \xmem_inst/mem[3][24] ) );
  DFF_X1 \xmem_inst/mem_reg[3][23]  ( .D(n4264), .CK(clk), .QN(
        \xmem_inst/mem[3][23] ) );
  DFF_X1 \xmem_inst/mem_reg[3][22]  ( .D(n4263), .CK(clk), .QN(
        \xmem_inst/mem[3][22] ) );
  DFF_X1 \xmem_inst/mem_reg[3][21]  ( .D(n4262), .CK(clk), .QN(
        \xmem_inst/mem[3][21] ) );
  DFF_X1 \xmem_inst/mem_reg[3][20]  ( .D(n4261), .CK(clk), .QN(
        \xmem_inst/mem[3][20] ) );
  DFF_X1 \xmem_inst/mem_reg[3][18]  ( .D(n4259), .CK(clk), .QN(
        \xmem_inst/mem[3][18] ) );
  DFF_X1 \xmem_inst/mem_reg[3][17]  ( .D(n4258), .CK(clk), .QN(
        \xmem_inst/mem[3][17] ) );
  DFF_X1 \xmem_inst/mem_reg[3][16]  ( .D(n4257), .CK(clk), .QN(
        \xmem_inst/mem[3][16] ) );
  DFF_X1 \xmem_inst/mem_reg[3][13]  ( .D(n4254), .CK(clk), .QN(
        \xmem_inst/mem[3][13] ) );
  DFF_X1 \xmem_inst/mem_reg[3][12]  ( .D(n4253), .CK(clk), .QN(
        \xmem_inst/mem[3][12] ) );
  DFF_X1 \xmem_inst/mem_reg[3][10]  ( .D(n4251), .CK(clk), .QN(
        \xmem_inst/mem[3][10] ) );
  DFF_X1 \xmem_inst/mem_reg[3][4]  ( .D(n4245), .CK(clk), .QN(
        \xmem_inst/mem[3][4] ) );
  DFF_X1 \xmem_inst/mem_reg[3][3]  ( .D(n4244), .CK(clk), .QN(
        \xmem_inst/mem[3][3] ) );
  DFF_X1 \xmem_inst/mem_reg[3][2]  ( .D(n4243), .CK(clk), .QN(
        \xmem_inst/mem[3][2] ) );
  DFF_X1 \xmem_inst/mem_reg[3][1]  ( .D(n4242), .CK(clk), .QN(
        \xmem_inst/mem[3][1] ) );
  DFF_X1 \xmem_inst/mem_reg[3][0]  ( .D(n4241), .CK(clk), .QN(
        \xmem_inst/mem[3][0] ) );
  DFF_X1 \xmem_inst/mem_reg[2][28]  ( .D(n4237), .CK(clk), .QN(
        \xmem_inst/mem[2][28] ) );
  DFF_X1 \xmem_inst/mem_reg[2][26]  ( .D(n4235), .CK(clk), .QN(
        \xmem_inst/mem[2][26] ) );
  DFF_X1 \xmem_inst/mem_reg[2][24]  ( .D(n4233), .CK(clk), .QN(
        \xmem_inst/mem[2][24] ) );
  DFF_X1 \xmem_inst/mem_reg[2][23]  ( .D(n4232), .CK(clk), .QN(
        \xmem_inst/mem[2][23] ) );
  DFF_X1 \xmem_inst/mem_reg[2][22]  ( .D(n4231), .CK(clk), .QN(
        \xmem_inst/mem[2][22] ) );
  DFF_X1 \xmem_inst/mem_reg[2][21]  ( .D(n4230), .CK(clk), .QN(
        \xmem_inst/mem[2][21] ) );
  DFF_X1 \xmem_inst/mem_reg[2][20]  ( .D(n4229), .CK(clk), .QN(
        \xmem_inst/mem[2][20] ) );
  DFF_X1 \xmem_inst/mem_reg[2][18]  ( .D(n4227), .CK(clk), .QN(
        \xmem_inst/mem[2][18] ) );
  DFF_X1 \xmem_inst/mem_reg[2][17]  ( .D(n4226), .CK(clk), .QN(
        \xmem_inst/mem[2][17] ) );
  DFF_X1 \xmem_inst/mem_reg[2][16]  ( .D(n4225), .CK(clk), .QN(
        \xmem_inst/mem[2][16] ) );
  DFF_X1 \xmem_inst/mem_reg[2][13]  ( .D(n4222), .CK(clk), .QN(
        \xmem_inst/mem[2][13] ) );
  DFF_X1 \xmem_inst/mem_reg[2][12]  ( .D(n4221), .CK(clk), .QN(
        \xmem_inst/mem[2][12] ) );
  DFF_X1 \xmem_inst/mem_reg[2][10]  ( .D(n4219), .CK(clk), .QN(
        \xmem_inst/mem[2][10] ) );
  DFF_X1 \xmem_inst/mem_reg[2][4]  ( .D(n4213), .CK(clk), .QN(
        \xmem_inst/mem[2][4] ) );
  DFF_X1 \xmem_inst/mem_reg[2][3]  ( .D(n4212), .CK(clk), .QN(
        \xmem_inst/mem[2][3] ) );
  DFF_X1 \xmem_inst/mem_reg[2][2]  ( .D(n4211), .CK(clk), .QN(
        \xmem_inst/mem[2][2] ) );
  DFF_X1 \xmem_inst/mem_reg[2][1]  ( .D(n4210), .CK(clk), .QN(
        \xmem_inst/mem[2][1] ) );
  DFF_X1 \xmem_inst/mem_reg[2][0]  ( .D(n4209), .CK(clk), .QN(
        \xmem_inst/mem[2][0] ) );
  DFF_X1 \xmem_inst/mem_reg[17][28]  ( .D(n4716), .CK(clk), .QN(
        \xmem_inst/mem[17][28] ) );
  DFF_X1 \xmem_inst/mem_reg[17][26]  ( .D(n4714), .CK(clk), .QN(
        \xmem_inst/mem[17][26] ) );
  DFF_X1 \xmem_inst/mem_reg[17][24]  ( .D(n4712), .CK(clk), .QN(
        \xmem_inst/mem[17][24] ) );
  DFF_X1 \xmem_inst/mem_reg[17][23]  ( .D(n4711), .CK(clk), .QN(
        \xmem_inst/mem[17][23] ) );
  DFF_X1 \xmem_inst/mem_reg[17][22]  ( .D(n4710), .CK(clk), .QN(
        \xmem_inst/mem[17][22] ) );
  DFF_X1 \xmem_inst/mem_reg[17][21]  ( .D(n4709), .CK(clk), .QN(
        \xmem_inst/mem[17][21] ) );
  DFF_X1 \xmem_inst/mem_reg[17][20]  ( .D(n4708), .CK(clk), .QN(
        \xmem_inst/mem[17][20] ) );
  DFF_X1 \xmem_inst/mem_reg[17][18]  ( .D(n4706), .CK(clk), .QN(
        \xmem_inst/mem[17][18] ) );
  DFF_X1 \xmem_inst/mem_reg[17][17]  ( .D(n4705), .CK(clk), .QN(
        \xmem_inst/mem[17][17] ) );
  DFF_X1 \xmem_inst/mem_reg[17][16]  ( .D(n4704), .CK(clk), .QN(
        \xmem_inst/mem[17][16] ) );
  DFF_X1 \xmem_inst/mem_reg[17][13]  ( .D(n4701), .CK(clk), .QN(
        \xmem_inst/mem[17][13] ) );
  DFF_X1 \xmem_inst/mem_reg[17][12]  ( .D(n4700), .CK(clk), .QN(
        \xmem_inst/mem[17][12] ) );
  DFF_X1 \xmem_inst/mem_reg[17][10]  ( .D(n4698), .CK(clk), .QN(
        \xmem_inst/mem[17][10] ) );
  DFF_X1 \xmem_inst/mem_reg[17][4]  ( .D(n4692), .CK(clk), .QN(
        \xmem_inst/mem[17][4] ) );
  DFF_X1 \xmem_inst/mem_reg[17][3]  ( .D(n4691), .CK(clk), .QN(
        \xmem_inst/mem[17][3] ) );
  DFF_X1 \xmem_inst/mem_reg[17][2]  ( .D(n4690), .CK(clk), .QN(
        \xmem_inst/mem[17][2] ) );
  DFF_X1 \xmem_inst/mem_reg[17][1]  ( .D(n4689), .CK(clk), .QN(
        \xmem_inst/mem[17][1] ) );
  DFF_X1 \xmem_inst/mem_reg[17][0]  ( .D(n4688), .CK(clk), .QN(
        \xmem_inst/mem[17][0] ) );
  DFF_X1 \xmem_inst/mem_reg[16][28]  ( .D(n4684), .CK(clk), .QN(
        \xmem_inst/mem[16][28] ) );
  DFF_X1 \xmem_inst/mem_reg[16][26]  ( .D(n4682), .CK(clk), .QN(
        \xmem_inst/mem[16][26] ) );
  DFF_X1 \xmem_inst/mem_reg[16][24]  ( .D(n4680), .CK(clk), .QN(
        \xmem_inst/mem[16][24] ) );
  DFF_X1 \xmem_inst/mem_reg[16][23]  ( .D(n4679), .CK(clk), .QN(
        \xmem_inst/mem[16][23] ) );
  DFF_X1 \xmem_inst/mem_reg[16][22]  ( .D(n4678), .CK(clk), .QN(
        \xmem_inst/mem[16][22] ) );
  DFF_X1 \xmem_inst/mem_reg[16][21]  ( .D(n4677), .CK(clk), .QN(
        \xmem_inst/mem[16][21] ) );
  DFF_X1 \xmem_inst/mem_reg[16][20]  ( .D(n4676), .CK(clk), .QN(
        \xmem_inst/mem[16][20] ) );
  DFF_X1 \xmem_inst/mem_reg[16][18]  ( .D(n4674), .CK(clk), .QN(
        \xmem_inst/mem[16][18] ) );
  DFF_X1 \xmem_inst/mem_reg[16][17]  ( .D(n4673), .CK(clk), .QN(
        \xmem_inst/mem[16][17] ) );
  DFF_X1 \xmem_inst/mem_reg[16][16]  ( .D(n4672), .CK(clk), .QN(
        \xmem_inst/mem[16][16] ) );
  DFF_X1 \xmem_inst/mem_reg[16][13]  ( .D(n4669), .CK(clk), .QN(
        \xmem_inst/mem[16][13] ) );
  DFF_X1 \xmem_inst/mem_reg[16][12]  ( .D(n4668), .CK(clk), .QN(
        \xmem_inst/mem[16][12] ) );
  DFF_X1 \xmem_inst/mem_reg[16][10]  ( .D(n4666), .CK(clk), .QN(
        \xmem_inst/mem[16][10] ) );
  DFF_X1 \xmem_inst/mem_reg[16][4]  ( .D(n4660), .CK(clk), .QN(
        \xmem_inst/mem[16][4] ) );
  DFF_X1 \xmem_inst/mem_reg[16][3]  ( .D(n4659), .CK(clk), .QN(
        \xmem_inst/mem[16][3] ) );
  DFF_X1 \xmem_inst/mem_reg[16][2]  ( .D(n4658), .CK(clk), .QN(
        \xmem_inst/mem[16][2] ) );
  DFF_X1 \xmem_inst/mem_reg[16][1]  ( .D(n4657), .CK(clk), .QN(
        \xmem_inst/mem[16][1] ) );
  DFF_X1 \xmem_inst/mem_reg[16][0]  ( .D(n4656), .CK(clk), .QN(
        \xmem_inst/mem[16][0] ) );
  DFF_X1 \xmem_inst/mem_reg[1][28]  ( .D(n4205), .CK(clk), .QN(
        \xmem_inst/mem[1][28] ) );
  DFF_X1 \xmem_inst/mem_reg[1][26]  ( .D(n4203), .CK(clk), .QN(
        \xmem_inst/mem[1][26] ) );
  DFF_X1 \xmem_inst/mem_reg[1][24]  ( .D(n4201), .CK(clk), .QN(
        \xmem_inst/mem[1][24] ) );
  DFF_X1 \xmem_inst/mem_reg[1][23]  ( .D(n4200), .CK(clk), .QN(
        \xmem_inst/mem[1][23] ) );
  DFF_X1 \xmem_inst/mem_reg[1][22]  ( .D(n4199), .CK(clk), .QN(
        \xmem_inst/mem[1][22] ) );
  DFF_X1 \xmem_inst/mem_reg[1][21]  ( .D(n4198), .CK(clk), .QN(
        \xmem_inst/mem[1][21] ) );
  DFF_X1 \xmem_inst/mem_reg[1][20]  ( .D(n4197), .CK(clk), .QN(
        \xmem_inst/mem[1][20] ) );
  DFF_X1 \xmem_inst/mem_reg[1][18]  ( .D(n4195), .CK(clk), .QN(
        \xmem_inst/mem[1][18] ) );
  DFF_X1 \xmem_inst/mem_reg[1][17]  ( .D(n4194), .CK(clk), .QN(
        \xmem_inst/mem[1][17] ) );
  DFF_X1 \xmem_inst/mem_reg[1][16]  ( .D(n4193), .CK(clk), .QN(
        \xmem_inst/mem[1][16] ) );
  DFF_X1 \xmem_inst/mem_reg[1][13]  ( .D(n4190), .CK(clk), .QN(
        \xmem_inst/mem[1][13] ) );
  DFF_X1 \xmem_inst/mem_reg[1][12]  ( .D(n4189), .CK(clk), .QN(
        \xmem_inst/mem[1][12] ) );
  DFF_X1 \xmem_inst/mem_reg[1][10]  ( .D(n4187), .CK(clk), .QN(
        \xmem_inst/mem[1][10] ) );
  DFF_X1 \xmem_inst/mem_reg[1][4]  ( .D(n4181), .CK(clk), .QN(
        \xmem_inst/mem[1][4] ) );
  DFF_X1 \xmem_inst/mem_reg[1][3]  ( .D(n4180), .CK(clk), .QN(
        \xmem_inst/mem[1][3] ) );
  DFF_X1 \xmem_inst/mem_reg[1][2]  ( .D(n4179), .CK(clk), .QN(
        \xmem_inst/mem[1][2] ) );
  DFF_X1 \xmem_inst/mem_reg[1][1]  ( .D(n4178), .CK(clk), .QN(
        \xmem_inst/mem[1][1] ) );
  DFF_X1 \xmem_inst/mem_reg[1][0]  ( .D(n4177), .CK(clk), .QN(
        \xmem_inst/mem[1][0] ) );
  DFF_X1 \xmem_inst/mem_reg[0][28]  ( .D(n4173), .CK(clk), .QN(
        \xmem_inst/mem[0][28] ) );
  DFF_X1 \xmem_inst/mem_reg[0][26]  ( .D(n4171), .CK(clk), .QN(
        \xmem_inst/mem[0][26] ) );
  DFF_X1 \xmem_inst/mem_reg[0][24]  ( .D(n4169), .CK(clk), .QN(
        \xmem_inst/mem[0][24] ) );
  DFF_X1 \xmem_inst/mem_reg[0][23]  ( .D(n4168), .CK(clk), .QN(
        \xmem_inst/mem[0][23] ) );
  DFF_X1 \xmem_inst/mem_reg[0][22]  ( .D(n4167), .CK(clk), .QN(
        \xmem_inst/mem[0][22] ) );
  DFF_X1 \xmem_inst/mem_reg[0][21]  ( .D(n4166), .CK(clk), .QN(
        \xmem_inst/mem[0][21] ) );
  DFF_X1 \xmem_inst/mem_reg[0][20]  ( .D(n4165), .CK(clk), .QN(
        \xmem_inst/mem[0][20] ) );
  DFF_X1 \xmem_inst/mem_reg[0][18]  ( .D(n4163), .CK(clk), .QN(
        \xmem_inst/mem[0][18] ) );
  DFF_X1 \xmem_inst/mem_reg[0][17]  ( .D(n4162), .CK(clk), .QN(
        \xmem_inst/mem[0][17] ) );
  DFF_X1 \xmem_inst/mem_reg[0][16]  ( .D(n4161), .CK(clk), .QN(
        \xmem_inst/mem[0][16] ) );
  DFF_X1 \xmem_inst/mem_reg[0][13]  ( .D(n4158), .CK(clk), .QN(
        \xmem_inst/mem[0][13] ) );
  DFF_X1 \xmem_inst/mem_reg[0][12]  ( .D(n4157), .CK(clk), .QN(
        \xmem_inst/mem[0][12] ) );
  DFF_X1 \xmem_inst/mem_reg[0][10]  ( .D(n4155), .CK(clk), .QN(
        \xmem_inst/mem[0][10] ) );
  DFF_X1 \xmem_inst/mem_reg[0][4]  ( .D(n4149), .CK(clk), .QN(
        \xmem_inst/mem[0][4] ) );
  DFF_X1 \xmem_inst/mem_reg[0][3]  ( .D(n4148), .CK(clk), .QN(
        \xmem_inst/mem[0][3] ) );
  DFF_X1 \xmem_inst/mem_reg[0][2]  ( .D(n4147), .CK(clk), .QN(
        \xmem_inst/mem[0][2] ) );
  DFF_X1 \xmem_inst/mem_reg[0][1]  ( .D(n4146), .CK(clk), .QN(
        \xmem_inst/mem[0][1] ) );
  DFF_X1 \xmem_inst/mem_reg[0][0]  ( .D(n4145), .CK(clk), .QN(
        \xmem_inst/mem[0][0] ) );
  DFF_X1 \xmem_inst/mem_reg[18][29]  ( .D(n4749), .CK(clk), .QN(
        \xmem_inst/mem[18][29] ) );
  DFF_X1 \xmem_inst/mem_reg[18][27]  ( .D(n4747), .CK(clk), .QN(
        \xmem_inst/mem[18][27] ) );
  DFF_X1 \xmem_inst/mem_reg[18][25]  ( .D(n4745), .CK(clk), .QN(
        \xmem_inst/mem[18][25] ) );
  DFF_X1 \xmem_inst/mem_reg[18][14]  ( .D(n4734), .CK(clk), .QN(
        \xmem_inst/mem[18][14] ) );
  DFF_X1 \xmem_inst/mem_reg[18][11]  ( .D(n4731), .CK(clk), .QN(
        \xmem_inst/mem[18][11] ) );
  DFF_X1 \xmem_inst/mem_reg[18][9]  ( .D(n4729), .CK(clk), .QN(
        \xmem_inst/mem[18][9] ) );
  DFF_X1 \xmem_inst/mem_reg[18][8]  ( .D(n4728), .CK(clk), .QN(
        \xmem_inst/mem[18][8] ) );
  DFF_X1 \xmem_inst/mem_reg[18][7]  ( .D(n4727), .CK(clk), .QN(
        \xmem_inst/mem[18][7] ) );
  DFF_X1 \xmem_inst/mem_reg[18][6]  ( .D(n4726), .CK(clk), .QN(
        \xmem_inst/mem[18][6] ) );
  DFF_X1 \xmem_inst/mem_reg[18][5]  ( .D(n4725), .CK(clk), .QN(
        \xmem_inst/mem[18][5] ) );
  DFF_X1 \xmem_inst/mem_reg[2][29]  ( .D(n4238), .CK(clk), .QN(
        \xmem_inst/mem[2][29] ) );
  DFF_X1 \xmem_inst/mem_reg[2][27]  ( .D(n4236), .CK(clk), .QN(
        \xmem_inst/mem[2][27] ) );
  DFF_X1 \xmem_inst/mem_reg[2][25]  ( .D(n4234), .CK(clk), .QN(
        \xmem_inst/mem[2][25] ) );
  DFF_X1 \xmem_inst/mem_reg[2][14]  ( .D(n4223), .CK(clk), .QN(
        \xmem_inst/mem[2][14] ) );
  DFF_X1 \xmem_inst/mem_reg[2][11]  ( .D(n4220), .CK(clk), .QN(
        \xmem_inst/mem[2][11] ) );
  DFF_X1 \xmem_inst/mem_reg[2][9]  ( .D(n4218), .CK(clk), .QN(
        \xmem_inst/mem[2][9] ) );
  DFF_X1 \xmem_inst/mem_reg[2][8]  ( .D(n4217), .CK(clk), .QN(
        \xmem_inst/mem[2][8] ) );
  DFF_X1 \xmem_inst/mem_reg[2][7]  ( .D(n4216), .CK(clk), .QN(
        \xmem_inst/mem[2][7] ) );
  DFF_X1 \xmem_inst/mem_reg[2][6]  ( .D(n4215), .CK(clk), .QN(
        \xmem_inst/mem[2][6] ) );
  DFF_X1 \xmem_inst/mem_reg[2][5]  ( .D(n4214), .CK(clk), .QN(
        \xmem_inst/mem[2][5] ) );
  DFF_X1 \xmem_inst/mem_reg[17][29]  ( .D(n4717), .CK(clk), .QN(
        \xmem_inst/mem[17][29] ) );
  DFF_X1 \xmem_inst/mem_reg[17][27]  ( .D(n4715), .CK(clk), .QN(
        \xmem_inst/mem[17][27] ) );
  DFF_X1 \xmem_inst/mem_reg[17][25]  ( .D(n4713), .CK(clk), .QN(
        \xmem_inst/mem[17][25] ) );
  DFF_X1 \xmem_inst/mem_reg[17][14]  ( .D(n4702), .CK(clk), .QN(
        \xmem_inst/mem[17][14] ) );
  DFF_X1 \xmem_inst/mem_reg[17][11]  ( .D(n4699), .CK(clk), .QN(
        \xmem_inst/mem[17][11] ) );
  DFF_X1 \xmem_inst/mem_reg[17][9]  ( .D(n4697), .CK(clk), .QN(
        \xmem_inst/mem[17][9] ) );
  DFF_X1 \xmem_inst/mem_reg[17][8]  ( .D(n4696), .CK(clk), .QN(
        \xmem_inst/mem[17][8] ) );
  DFF_X1 \xmem_inst/mem_reg[17][7]  ( .D(n4695), .CK(clk), .QN(
        \xmem_inst/mem[17][7] ) );
  DFF_X1 \xmem_inst/mem_reg[17][6]  ( .D(n4694), .CK(clk), .QN(
        \xmem_inst/mem[17][6] ) );
  DFF_X1 \xmem_inst/mem_reg[17][5]  ( .D(n4693), .CK(clk), .QN(
        \xmem_inst/mem[17][5] ) );
  DFF_X1 \xmem_inst/mem_reg[16][29]  ( .D(n4685), .CK(clk), .QN(
        \xmem_inst/mem[16][29] ) );
  DFF_X1 \xmem_inst/mem_reg[16][27]  ( .D(n4683), .CK(clk), .QN(
        \xmem_inst/mem[16][27] ) );
  DFF_X1 \xmem_inst/mem_reg[16][25]  ( .D(n4681), .CK(clk), .QN(
        \xmem_inst/mem[16][25] ) );
  DFF_X1 \xmem_inst/mem_reg[16][14]  ( .D(n4670), .CK(clk), .QN(
        \xmem_inst/mem[16][14] ) );
  DFF_X1 \xmem_inst/mem_reg[16][11]  ( .D(n4667), .CK(clk), .QN(
        \xmem_inst/mem[16][11] ) );
  DFF_X1 \xmem_inst/mem_reg[16][9]  ( .D(n4665), .CK(clk), .QN(
        \xmem_inst/mem[16][9] ) );
  DFF_X1 \xmem_inst/mem_reg[16][8]  ( .D(n4664), .CK(clk), .QN(
        \xmem_inst/mem[16][8] ) );
  DFF_X1 \xmem_inst/mem_reg[16][7]  ( .D(n4663), .CK(clk), .QN(
        \xmem_inst/mem[16][7] ) );
  DFF_X1 \xmem_inst/mem_reg[16][6]  ( .D(n4662), .CK(clk), .QN(
        \xmem_inst/mem[16][6] ) );
  DFF_X1 \xmem_inst/mem_reg[16][5]  ( .D(n4661), .CK(clk), .QN(
        \xmem_inst/mem[16][5] ) );
  DFF_X1 \xmem_inst/mem_reg[1][29]  ( .D(n4206), .CK(clk), .QN(
        \xmem_inst/mem[1][29] ) );
  DFF_X1 \xmem_inst/mem_reg[1][27]  ( .D(n4204), .CK(clk), .QN(
        \xmem_inst/mem[1][27] ) );
  DFF_X1 \xmem_inst/mem_reg[1][25]  ( .D(n4202), .CK(clk), .QN(
        \xmem_inst/mem[1][25] ) );
  DFF_X1 \xmem_inst/mem_reg[1][14]  ( .D(n4191), .CK(clk), .QN(
        \xmem_inst/mem[1][14] ) );
  DFF_X1 \xmem_inst/mem_reg[1][11]  ( .D(n4188), .CK(clk), .QN(
        \xmem_inst/mem[1][11] ) );
  DFF_X1 \xmem_inst/mem_reg[1][9]  ( .D(n4186), .CK(clk), .QN(
        \xmem_inst/mem[1][9] ) );
  DFF_X1 \xmem_inst/mem_reg[1][8]  ( .D(n4185), .CK(clk), .QN(
        \xmem_inst/mem[1][8] ) );
  DFF_X1 \xmem_inst/mem_reg[1][7]  ( .D(n4184), .CK(clk), .QN(
        \xmem_inst/mem[1][7] ) );
  DFF_X1 \xmem_inst/mem_reg[1][6]  ( .D(n4183), .CK(clk), .QN(
        \xmem_inst/mem[1][6] ) );
  DFF_X1 \xmem_inst/mem_reg[1][5]  ( .D(n4182), .CK(clk), .QN(
        \xmem_inst/mem[1][5] ) );
  DFF_X1 \xmem_inst/mem_reg[0][29]  ( .D(n4174), .CK(clk), .QN(
        \xmem_inst/mem[0][29] ) );
  DFF_X1 \xmem_inst/mem_reg[0][27]  ( .D(n4172), .CK(clk), .QN(
        \xmem_inst/mem[0][27] ) );
  DFF_X1 \xmem_inst/mem_reg[0][25]  ( .D(n4170), .CK(clk), .QN(
        \xmem_inst/mem[0][25] ) );
  DFF_X1 \xmem_inst/mem_reg[0][14]  ( .D(n4159), .CK(clk), .QN(
        \xmem_inst/mem[0][14] ) );
  DFF_X1 \xmem_inst/mem_reg[0][11]  ( .D(n4156), .CK(clk), .QN(
        \xmem_inst/mem[0][11] ) );
  DFF_X1 \xmem_inst/mem_reg[0][9]  ( .D(n4154), .CK(clk), .QN(
        \xmem_inst/mem[0][9] ) );
  DFF_X1 \xmem_inst/mem_reg[0][8]  ( .D(n4153), .CK(clk), .QN(
        \xmem_inst/mem[0][8] ) );
  DFF_X1 \xmem_inst/mem_reg[0][7]  ( .D(n4152), .CK(clk), .QN(
        \xmem_inst/mem[0][7] ) );
  DFF_X1 \xmem_inst/mem_reg[0][6]  ( .D(n4151), .CK(clk), .QN(
        \xmem_inst/mem[0][6] ) );
  DFF_X1 \xmem_inst/mem_reg[0][5]  ( .D(n4150), .CK(clk), .QN(
        \xmem_inst/mem[0][5] ) );
  DFF_X1 \xmem_inst/mem_reg[31][31]  ( .D(n5167), .CK(clk), .QN(
        \xmem_inst/mem[31][31] ) );
  DFF_X1 \xmem_inst/mem_reg[31][30]  ( .D(n5166), .CK(clk), .QN(
        \xmem_inst/mem[31][30] ) );
  DFF_X1 \xmem_inst/mem_reg[31][19]  ( .D(n5155), .CK(clk), .QN(
        \xmem_inst/mem[31][19] ) );
  DFF_X1 \xmem_inst/mem_reg[31][15]  ( .D(n5151), .CK(clk), .QN(
        \xmem_inst/mem[31][15] ) );
  DFF_X1 \xmem_inst/mem_reg[15][31]  ( .D(n4655), .CK(clk), .QN(
        \xmem_inst/mem[15][31] ) );
  DFF_X1 \xmem_inst/mem_reg[15][30]  ( .D(n4654), .CK(clk), .QN(
        \xmem_inst/mem[15][30] ) );
  DFF_X1 \xmem_inst/mem_reg[15][19]  ( .D(n4643), .CK(clk), .QN(
        \xmem_inst/mem[15][19] ) );
  DFF_X1 \xmem_inst/mem_reg[15][15]  ( .D(n4639), .CK(clk), .QN(
        \xmem_inst/mem[15][15] ) );
  DFF_X1 \xmem_inst/mem_reg[27][31]  ( .D(n5039), .CK(clk), .QN(
        \xmem_inst/mem[27][31] ) );
  DFF_X1 \xmem_inst/mem_reg[27][30]  ( .D(n5038), .CK(clk), .QN(
        \xmem_inst/mem[27][30] ) );
  DFF_X1 \xmem_inst/mem_reg[27][19]  ( .D(n5027), .CK(clk), .QN(
        \xmem_inst/mem[27][19] ) );
  DFF_X1 \xmem_inst/mem_reg[27][15]  ( .D(n5023), .CK(clk), .QN(
        \xmem_inst/mem[27][15] ) );
  DFF_X1 \xmem_inst/mem_reg[11][31]  ( .D(n4527), .CK(clk), .QN(
        \xmem_inst/mem[11][31] ) );
  DFF_X1 \xmem_inst/mem_reg[11][30]  ( .D(n4526), .CK(clk), .QN(
        \xmem_inst/mem[11][30] ) );
  DFF_X1 \xmem_inst/mem_reg[11][19]  ( .D(n4515), .CK(clk), .QN(
        \xmem_inst/mem[11][19] ) );
  DFF_X1 \xmem_inst/mem_reg[11][15]  ( .D(n4511), .CK(clk), .QN(
        \xmem_inst/mem[11][15] ) );
  DFF_X1 \xmem_inst/mem_reg[30][31]  ( .D(n5135), .CK(clk), .QN(
        \xmem_inst/mem[30][31] ) );
  DFF_X1 \xmem_inst/mem_reg[30][30]  ( .D(n5134), .CK(clk), .QN(
        \xmem_inst/mem[30][30] ) );
  DFF_X1 \xmem_inst/mem_reg[30][19]  ( .D(n5123), .CK(clk), .QN(
        \xmem_inst/mem[30][19] ) );
  DFF_X1 \xmem_inst/mem_reg[30][15]  ( .D(n5119), .CK(clk), .QN(
        \xmem_inst/mem[30][15] ) );
  DFF_X1 \xmem_inst/mem_reg[29][31]  ( .D(n5103), .CK(clk), .QN(
        \xmem_inst/mem[29][31] ) );
  DFF_X1 \xmem_inst/mem_reg[29][30]  ( .D(n5102), .CK(clk), .QN(
        \xmem_inst/mem[29][30] ) );
  DFF_X1 \xmem_inst/mem_reg[29][19]  ( .D(n5091), .CK(clk), .QN(
        \xmem_inst/mem[29][19] ) );
  DFF_X1 \xmem_inst/mem_reg[29][15]  ( .D(n5087), .CK(clk), .QN(
        \xmem_inst/mem[29][15] ) );
  DFF_X1 \xmem_inst/mem_reg[28][31]  ( .D(n5071), .CK(clk), .QN(
        \xmem_inst/mem[28][31] ) );
  DFF_X1 \xmem_inst/mem_reg[28][30]  ( .D(n5070), .CK(clk), .QN(
        \xmem_inst/mem[28][30] ) );
  DFF_X1 \xmem_inst/mem_reg[28][19]  ( .D(n5059), .CK(clk), .QN(
        \xmem_inst/mem[28][19] ) );
  DFF_X1 \xmem_inst/mem_reg[28][15]  ( .D(n5055), .CK(clk), .QN(
        \xmem_inst/mem[28][15] ) );
  DFF_X1 \xmem_inst/mem_reg[14][31]  ( .D(n4623), .CK(clk), .QN(
        \xmem_inst/mem[14][31] ) );
  DFF_X1 \xmem_inst/mem_reg[14][30]  ( .D(n4622), .CK(clk), .QN(
        \xmem_inst/mem[14][30] ) );
  DFF_X1 \xmem_inst/mem_reg[14][19]  ( .D(n4611), .CK(clk), .QN(
        \xmem_inst/mem[14][19] ) );
  DFF_X1 \xmem_inst/mem_reg[14][15]  ( .D(n4607), .CK(clk), .QN(
        \xmem_inst/mem[14][15] ) );
  DFF_X1 \xmem_inst/mem_reg[13][31]  ( .D(n4591), .CK(clk), .QN(
        \xmem_inst/mem[13][31] ) );
  DFF_X1 \xmem_inst/mem_reg[13][30]  ( .D(n4590), .CK(clk), .QN(
        \xmem_inst/mem[13][30] ) );
  DFF_X1 \xmem_inst/mem_reg[13][19]  ( .D(n4579), .CK(clk), .QN(
        \xmem_inst/mem[13][19] ) );
  DFF_X1 \xmem_inst/mem_reg[13][15]  ( .D(n4575), .CK(clk), .QN(
        \xmem_inst/mem[13][15] ) );
  DFF_X1 \xmem_inst/mem_reg[12][31]  ( .D(n4559), .CK(clk), .QN(
        \xmem_inst/mem[12][31] ) );
  DFF_X1 \xmem_inst/mem_reg[12][30]  ( .D(n4558), .CK(clk), .QN(
        \xmem_inst/mem[12][30] ) );
  DFF_X1 \xmem_inst/mem_reg[12][19]  ( .D(n4547), .CK(clk), .QN(
        \xmem_inst/mem[12][19] ) );
  DFF_X1 \xmem_inst/mem_reg[12][15]  ( .D(n4543), .CK(clk), .QN(
        \xmem_inst/mem[12][15] ) );
  DFF_X1 \xmem_inst/mem_reg[26][31]  ( .D(n5007), .CK(clk), .QN(
        \xmem_inst/mem[26][31] ) );
  DFF_X1 \xmem_inst/mem_reg[26][30]  ( .D(n5006), .CK(clk), .QN(
        \xmem_inst/mem[26][30] ) );
  DFF_X1 \xmem_inst/mem_reg[26][19]  ( .D(n4995), .CK(clk), .QN(
        \xmem_inst/mem[26][19] ) );
  DFF_X1 \xmem_inst/mem_reg[26][15]  ( .D(n4991), .CK(clk), .QN(
        \xmem_inst/mem[26][15] ) );
  DFF_X1 \xmem_inst/mem_reg[25][31]  ( .D(n4975), .CK(clk), .QN(
        \xmem_inst/mem[25][31] ) );
  DFF_X1 \xmem_inst/mem_reg[25][30]  ( .D(n4974), .CK(clk), .QN(
        \xmem_inst/mem[25][30] ) );
  DFF_X1 \xmem_inst/mem_reg[25][19]  ( .D(n4963), .CK(clk), .QN(
        \xmem_inst/mem[25][19] ) );
  DFF_X1 \xmem_inst/mem_reg[25][15]  ( .D(n4959), .CK(clk), .QN(
        \xmem_inst/mem[25][15] ) );
  DFF_X1 \xmem_inst/mem_reg[24][31]  ( .D(n4943), .CK(clk), .QN(
        \xmem_inst/mem[24][31] ) );
  DFF_X1 \xmem_inst/mem_reg[24][30]  ( .D(n4942), .CK(clk), .QN(
        \xmem_inst/mem[24][30] ) );
  DFF_X1 \xmem_inst/mem_reg[24][19]  ( .D(n4931), .CK(clk), .QN(
        \xmem_inst/mem[24][19] ) );
  DFF_X1 \xmem_inst/mem_reg[24][15]  ( .D(n4927), .CK(clk), .QN(
        \xmem_inst/mem[24][15] ) );
  DFF_X1 \xmem_inst/mem_reg[10][31]  ( .D(n4495), .CK(clk), .QN(
        \xmem_inst/mem[10][31] ) );
  DFF_X1 \xmem_inst/mem_reg[10][30]  ( .D(n4494), .CK(clk), .QN(
        \xmem_inst/mem[10][30] ) );
  DFF_X1 \xmem_inst/mem_reg[10][19]  ( .D(n4483), .CK(clk), .QN(
        \xmem_inst/mem[10][19] ) );
  DFF_X1 \xmem_inst/mem_reg[10][15]  ( .D(n4479), .CK(clk), .QN(
        \xmem_inst/mem[10][15] ) );
  DFF_X1 \xmem_inst/mem_reg[9][31]  ( .D(n4463), .CK(clk), .QN(
        \xmem_inst/mem[9][31] ) );
  DFF_X1 \xmem_inst/mem_reg[9][30]  ( .D(n4462), .CK(clk), .QN(
        \xmem_inst/mem[9][30] ) );
  DFF_X1 \xmem_inst/mem_reg[9][19]  ( .D(n4451), .CK(clk), .QN(
        \xmem_inst/mem[9][19] ) );
  DFF_X1 \xmem_inst/mem_reg[9][15]  ( .D(n4447), .CK(clk), .QN(
        \xmem_inst/mem[9][15] ) );
  DFF_X1 \xmem_inst/mem_reg[8][31]  ( .D(n4431), .CK(clk), .QN(
        \xmem_inst/mem[8][31] ) );
  DFF_X1 \xmem_inst/mem_reg[8][30]  ( .D(n4430), .CK(clk), .QN(
        \xmem_inst/mem[8][30] ) );
  DFF_X1 \xmem_inst/mem_reg[8][19]  ( .D(n4419), .CK(clk), .QN(
        \xmem_inst/mem[8][19] ) );
  DFF_X1 \xmem_inst/mem_reg[8][15]  ( .D(n4415), .CK(clk), .QN(
        \xmem_inst/mem[8][15] ) );
  DFF_X1 \xmem_inst/mem_reg[31][29]  ( .D(n5165), .CK(clk), .QN(
        \xmem_inst/mem[31][29] ) );
  DFF_X1 \xmem_inst/mem_reg[31][27]  ( .D(n5163), .CK(clk), .QN(
        \xmem_inst/mem[31][27] ) );
  DFF_X1 \xmem_inst/mem_reg[31][25]  ( .D(n5161), .CK(clk), .QN(
        \xmem_inst/mem[31][25] ) );
  DFF_X1 \xmem_inst/mem_reg[31][14]  ( .D(n5150), .CK(clk), .QN(
        \xmem_inst/mem[31][14] ) );
  DFF_X1 \xmem_inst/mem_reg[31][11]  ( .D(n5147), .CK(clk), .QN(
        \xmem_inst/mem[31][11] ) );
  DFF_X1 \xmem_inst/mem_reg[31][9]  ( .D(n5145), .CK(clk), .QN(
        \xmem_inst/mem[31][9] ) );
  DFF_X1 \xmem_inst/mem_reg[31][8]  ( .D(n5144), .CK(clk), .QN(
        \xmem_inst/mem[31][8] ) );
  DFF_X1 \xmem_inst/mem_reg[31][7]  ( .D(n5143), .CK(clk), .QN(
        \xmem_inst/mem[31][7] ) );
  DFF_X1 \xmem_inst/mem_reg[31][6]  ( .D(n5142), .CK(clk), .QN(
        \xmem_inst/mem[31][6] ) );
  DFF_X1 \xmem_inst/mem_reg[31][5]  ( .D(n5141), .CK(clk), .QN(
        \xmem_inst/mem[31][5] ) );
  DFF_X1 \xmem_inst/mem_reg[15][29]  ( .D(n4653), .CK(clk), .QN(
        \xmem_inst/mem[15][29] ) );
  DFF_X1 \xmem_inst/mem_reg[15][27]  ( .D(n4651), .CK(clk), .QN(
        \xmem_inst/mem[15][27] ) );
  DFF_X1 \xmem_inst/mem_reg[15][25]  ( .D(n4649), .CK(clk), .QN(
        \xmem_inst/mem[15][25] ) );
  DFF_X1 \xmem_inst/mem_reg[15][14]  ( .D(n4638), .CK(clk), .QN(
        \xmem_inst/mem[15][14] ) );
  DFF_X1 \xmem_inst/mem_reg[15][11]  ( .D(n4635), .CK(clk), .QN(
        \xmem_inst/mem[15][11] ) );
  DFF_X1 \xmem_inst/mem_reg[15][9]  ( .D(n4633), .CK(clk), .QN(
        \xmem_inst/mem[15][9] ) );
  DFF_X1 \xmem_inst/mem_reg[15][8]  ( .D(n4632), .CK(clk), .QN(
        \xmem_inst/mem[15][8] ) );
  DFF_X1 \xmem_inst/mem_reg[15][7]  ( .D(n4631), .CK(clk), .QN(
        \xmem_inst/mem[15][7] ) );
  DFF_X1 \xmem_inst/mem_reg[15][6]  ( .D(n4630), .CK(clk), .QN(
        \xmem_inst/mem[15][6] ) );
  DFF_X1 \xmem_inst/mem_reg[15][5]  ( .D(n4629), .CK(clk), .QN(
        \xmem_inst/mem[15][5] ) );
  DFF_X1 \xmem_inst/mem_reg[27][29]  ( .D(n5037), .CK(clk), .QN(
        \xmem_inst/mem[27][29] ) );
  DFF_X1 \xmem_inst/mem_reg[27][27]  ( .D(n5035), .CK(clk), .QN(
        \xmem_inst/mem[27][27] ) );
  DFF_X1 \xmem_inst/mem_reg[27][25]  ( .D(n5033), .CK(clk), .QN(
        \xmem_inst/mem[27][25] ) );
  DFF_X1 \xmem_inst/mem_reg[27][14]  ( .D(n5022), .CK(clk), .QN(
        \xmem_inst/mem[27][14] ) );
  DFF_X1 \xmem_inst/mem_reg[27][11]  ( .D(n5019), .CK(clk), .QN(
        \xmem_inst/mem[27][11] ) );
  DFF_X1 \xmem_inst/mem_reg[27][9]  ( .D(n5017), .CK(clk), .QN(
        \xmem_inst/mem[27][9] ) );
  DFF_X1 \xmem_inst/mem_reg[27][8]  ( .D(n5016), .CK(clk), .QN(
        \xmem_inst/mem[27][8] ) );
  DFF_X1 \xmem_inst/mem_reg[27][7]  ( .D(n5015), .CK(clk), .QN(
        \xmem_inst/mem[27][7] ) );
  DFF_X1 \xmem_inst/mem_reg[27][6]  ( .D(n5014), .CK(clk), .QN(
        \xmem_inst/mem[27][6] ) );
  DFF_X1 \xmem_inst/mem_reg[27][5]  ( .D(n5013), .CK(clk), .QN(
        \xmem_inst/mem[27][5] ) );
  DFF_X1 \xmem_inst/mem_reg[11][29]  ( .D(n4525), .CK(clk), .QN(
        \xmem_inst/mem[11][29] ) );
  DFF_X1 \xmem_inst/mem_reg[11][27]  ( .D(n4523), .CK(clk), .QN(
        \xmem_inst/mem[11][27] ) );
  DFF_X1 \xmem_inst/mem_reg[11][25]  ( .D(n4521), .CK(clk), .QN(
        \xmem_inst/mem[11][25] ) );
  DFF_X1 \xmem_inst/mem_reg[11][14]  ( .D(n4510), .CK(clk), .QN(
        \xmem_inst/mem[11][14] ) );
  DFF_X1 \xmem_inst/mem_reg[11][11]  ( .D(n4507), .CK(clk), .QN(
        \xmem_inst/mem[11][11] ) );
  DFF_X1 \xmem_inst/mem_reg[11][9]  ( .D(n4505), .CK(clk), .QN(
        \xmem_inst/mem[11][9] ) );
  DFF_X1 \xmem_inst/mem_reg[11][8]  ( .D(n4504), .CK(clk), .QN(
        \xmem_inst/mem[11][8] ) );
  DFF_X1 \xmem_inst/mem_reg[11][7]  ( .D(n4503), .CK(clk), .QN(
        \xmem_inst/mem[11][7] ) );
  DFF_X1 \xmem_inst/mem_reg[11][6]  ( .D(n4502), .CK(clk), .QN(
        \xmem_inst/mem[11][6] ) );
  DFF_X1 \xmem_inst/mem_reg[11][5]  ( .D(n4501), .CK(clk), .QN(
        \xmem_inst/mem[11][5] ) );
  DFF_X1 \xmem_inst/mem_reg[30][29]  ( .D(n5133), .CK(clk), .QN(
        \xmem_inst/mem[30][29] ) );
  DFF_X1 \xmem_inst/mem_reg[30][27]  ( .D(n5131), .CK(clk), .QN(
        \xmem_inst/mem[30][27] ) );
  DFF_X1 \xmem_inst/mem_reg[30][25]  ( .D(n5129), .CK(clk), .QN(
        \xmem_inst/mem[30][25] ) );
  DFF_X1 \xmem_inst/mem_reg[30][14]  ( .D(n5118), .CK(clk), .QN(
        \xmem_inst/mem[30][14] ) );
  DFF_X1 \xmem_inst/mem_reg[30][11]  ( .D(n5115), .CK(clk), .QN(
        \xmem_inst/mem[30][11] ) );
  DFF_X1 \xmem_inst/mem_reg[30][9]  ( .D(n5113), .CK(clk), .QN(
        \xmem_inst/mem[30][9] ) );
  DFF_X1 \xmem_inst/mem_reg[30][8]  ( .D(n5112), .CK(clk), .QN(
        \xmem_inst/mem[30][8] ) );
  DFF_X1 \xmem_inst/mem_reg[30][7]  ( .D(n5111), .CK(clk), .QN(
        \xmem_inst/mem[30][7] ) );
  DFF_X1 \xmem_inst/mem_reg[30][6]  ( .D(n5110), .CK(clk), .QN(
        \xmem_inst/mem[30][6] ) );
  DFF_X1 \xmem_inst/mem_reg[30][5]  ( .D(n5109), .CK(clk), .QN(
        \xmem_inst/mem[30][5] ) );
  DFF_X1 \xmem_inst/mem_reg[29][29]  ( .D(n5101), .CK(clk), .QN(
        \xmem_inst/mem[29][29] ) );
  DFF_X1 \xmem_inst/mem_reg[29][27]  ( .D(n5099), .CK(clk), .QN(
        \xmem_inst/mem[29][27] ) );
  DFF_X1 \xmem_inst/mem_reg[29][25]  ( .D(n5097), .CK(clk), .QN(
        \xmem_inst/mem[29][25] ) );
  DFF_X1 \xmem_inst/mem_reg[29][14]  ( .D(n5086), .CK(clk), .QN(
        \xmem_inst/mem[29][14] ) );
  DFF_X1 \xmem_inst/mem_reg[29][11]  ( .D(n5083), .CK(clk), .QN(
        \xmem_inst/mem[29][11] ) );
  DFF_X1 \xmem_inst/mem_reg[29][9]  ( .D(n5081), .CK(clk), .QN(
        \xmem_inst/mem[29][9] ) );
  DFF_X1 \xmem_inst/mem_reg[29][8]  ( .D(n5080), .CK(clk), .QN(
        \xmem_inst/mem[29][8] ) );
  DFF_X1 \xmem_inst/mem_reg[29][7]  ( .D(n5079), .CK(clk), .QN(
        \xmem_inst/mem[29][7] ) );
  DFF_X1 \xmem_inst/mem_reg[29][6]  ( .D(n5078), .CK(clk), .QN(
        \xmem_inst/mem[29][6] ) );
  DFF_X1 \xmem_inst/mem_reg[29][5]  ( .D(n5077), .CK(clk), .QN(
        \xmem_inst/mem[29][5] ) );
  DFF_X1 \xmem_inst/mem_reg[28][29]  ( .D(n5069), .CK(clk), .QN(
        \xmem_inst/mem[28][29] ) );
  DFF_X1 \xmem_inst/mem_reg[28][27]  ( .D(n5067), .CK(clk), .QN(
        \xmem_inst/mem[28][27] ) );
  DFF_X1 \xmem_inst/mem_reg[28][25]  ( .D(n5065), .CK(clk), .QN(
        \xmem_inst/mem[28][25] ) );
  DFF_X1 \xmem_inst/mem_reg[28][14]  ( .D(n5054), .CK(clk), .QN(
        \xmem_inst/mem[28][14] ) );
  DFF_X1 \xmem_inst/mem_reg[28][11]  ( .D(n5051), .CK(clk), .QN(
        \xmem_inst/mem[28][11] ) );
  DFF_X1 \xmem_inst/mem_reg[28][9]  ( .D(n5049), .CK(clk), .QN(
        \xmem_inst/mem[28][9] ) );
  DFF_X1 \xmem_inst/mem_reg[28][8]  ( .D(n5048), .CK(clk), .QN(
        \xmem_inst/mem[28][8] ) );
  DFF_X1 \xmem_inst/mem_reg[28][7]  ( .D(n5047), .CK(clk), .QN(
        \xmem_inst/mem[28][7] ) );
  DFF_X1 \xmem_inst/mem_reg[28][6]  ( .D(n5046), .CK(clk), .QN(
        \xmem_inst/mem[28][6] ) );
  DFF_X1 \xmem_inst/mem_reg[28][5]  ( .D(n5045), .CK(clk), .QN(
        \xmem_inst/mem[28][5] ) );
  DFF_X1 \xmem_inst/mem_reg[14][29]  ( .D(n4621), .CK(clk), .QN(
        \xmem_inst/mem[14][29] ) );
  DFF_X1 \xmem_inst/mem_reg[14][27]  ( .D(n4619), .CK(clk), .QN(
        \xmem_inst/mem[14][27] ) );
  DFF_X1 \xmem_inst/mem_reg[14][25]  ( .D(n4617), .CK(clk), .QN(
        \xmem_inst/mem[14][25] ) );
  DFF_X1 \xmem_inst/mem_reg[14][14]  ( .D(n4606), .CK(clk), .QN(
        \xmem_inst/mem[14][14] ) );
  DFF_X1 \xmem_inst/mem_reg[14][11]  ( .D(n4603), .CK(clk), .QN(
        \xmem_inst/mem[14][11] ) );
  DFF_X1 \xmem_inst/mem_reg[14][9]  ( .D(n4601), .CK(clk), .QN(
        \xmem_inst/mem[14][9] ) );
  DFF_X1 \xmem_inst/mem_reg[14][8]  ( .D(n4600), .CK(clk), .QN(
        \xmem_inst/mem[14][8] ) );
  DFF_X1 \xmem_inst/mem_reg[14][7]  ( .D(n4599), .CK(clk), .QN(
        \xmem_inst/mem[14][7] ) );
  DFF_X1 \xmem_inst/mem_reg[14][6]  ( .D(n4598), .CK(clk), .QN(
        \xmem_inst/mem[14][6] ) );
  DFF_X1 \xmem_inst/mem_reg[14][5]  ( .D(n4597), .CK(clk), .QN(
        \xmem_inst/mem[14][5] ) );
  DFF_X1 \xmem_inst/mem_reg[13][29]  ( .D(n4589), .CK(clk), .QN(
        \xmem_inst/mem[13][29] ) );
  DFF_X1 \xmem_inst/mem_reg[13][27]  ( .D(n4587), .CK(clk), .QN(
        \xmem_inst/mem[13][27] ) );
  DFF_X1 \xmem_inst/mem_reg[13][25]  ( .D(n4585), .CK(clk), .QN(
        \xmem_inst/mem[13][25] ) );
  DFF_X1 \xmem_inst/mem_reg[13][14]  ( .D(n4574), .CK(clk), .QN(
        \xmem_inst/mem[13][14] ) );
  DFF_X1 \xmem_inst/mem_reg[13][11]  ( .D(n4571), .CK(clk), .QN(
        \xmem_inst/mem[13][11] ) );
  DFF_X1 \xmem_inst/mem_reg[13][9]  ( .D(n4569), .CK(clk), .QN(
        \xmem_inst/mem[13][9] ) );
  DFF_X1 \xmem_inst/mem_reg[13][8]  ( .D(n4568), .CK(clk), .QN(
        \xmem_inst/mem[13][8] ) );
  DFF_X1 \xmem_inst/mem_reg[13][7]  ( .D(n4567), .CK(clk), .QN(
        \xmem_inst/mem[13][7] ) );
  DFF_X1 \xmem_inst/mem_reg[13][6]  ( .D(n4566), .CK(clk), .QN(
        \xmem_inst/mem[13][6] ) );
  DFF_X1 \xmem_inst/mem_reg[13][5]  ( .D(n4565), .CK(clk), .QN(
        \xmem_inst/mem[13][5] ) );
  DFF_X1 \xmem_inst/mem_reg[12][29]  ( .D(n4557), .CK(clk), .QN(
        \xmem_inst/mem[12][29] ) );
  DFF_X1 \xmem_inst/mem_reg[12][27]  ( .D(n4555), .CK(clk), .QN(
        \xmem_inst/mem[12][27] ) );
  DFF_X1 \xmem_inst/mem_reg[12][25]  ( .D(n4553), .CK(clk), .QN(
        \xmem_inst/mem[12][25] ) );
  DFF_X1 \xmem_inst/mem_reg[12][14]  ( .D(n4542), .CK(clk), .QN(
        \xmem_inst/mem[12][14] ) );
  DFF_X1 \xmem_inst/mem_reg[12][11]  ( .D(n4539), .CK(clk), .QN(
        \xmem_inst/mem[12][11] ) );
  DFF_X1 \xmem_inst/mem_reg[12][9]  ( .D(n4537), .CK(clk), .QN(
        \xmem_inst/mem[12][9] ) );
  DFF_X1 \xmem_inst/mem_reg[12][8]  ( .D(n4536), .CK(clk), .QN(
        \xmem_inst/mem[12][8] ) );
  DFF_X1 \xmem_inst/mem_reg[12][7]  ( .D(n4535), .CK(clk), .QN(
        \xmem_inst/mem[12][7] ) );
  DFF_X1 \xmem_inst/mem_reg[12][6]  ( .D(n4534), .CK(clk), .QN(
        \xmem_inst/mem[12][6] ) );
  DFF_X1 \xmem_inst/mem_reg[12][5]  ( .D(n4533), .CK(clk), .QN(
        \xmem_inst/mem[12][5] ) );
  DFF_X1 \xmem_inst/mem_reg[31][28]  ( .D(n5164), .CK(clk), .QN(
        \xmem_inst/mem[31][28] ) );
  DFF_X1 \xmem_inst/mem_reg[31][26]  ( .D(n5162), .CK(clk), .QN(
        \xmem_inst/mem[31][26] ) );
  DFF_X1 \xmem_inst/mem_reg[31][24]  ( .D(n5160), .CK(clk), .QN(
        \xmem_inst/mem[31][24] ) );
  DFF_X1 \xmem_inst/mem_reg[31][23]  ( .D(n5159), .CK(clk), .QN(
        \xmem_inst/mem[31][23] ) );
  DFF_X1 \xmem_inst/mem_reg[31][22]  ( .D(n5158), .CK(clk), .QN(
        \xmem_inst/mem[31][22] ) );
  DFF_X1 \xmem_inst/mem_reg[31][21]  ( .D(n5157), .CK(clk), .QN(
        \xmem_inst/mem[31][21] ) );
  DFF_X1 \xmem_inst/mem_reg[31][20]  ( .D(n5156), .CK(clk), .QN(
        \xmem_inst/mem[31][20] ) );
  DFF_X1 \xmem_inst/mem_reg[31][18]  ( .D(n5154), .CK(clk), .QN(
        \xmem_inst/mem[31][18] ) );
  DFF_X1 \xmem_inst/mem_reg[31][17]  ( .D(n5153), .CK(clk), .QN(
        \xmem_inst/mem[31][17] ) );
  DFF_X1 \xmem_inst/mem_reg[31][16]  ( .D(n5152), .CK(clk), .QN(
        \xmem_inst/mem[31][16] ) );
  DFF_X1 \xmem_inst/mem_reg[31][13]  ( .D(n5149), .CK(clk), .QN(
        \xmem_inst/mem[31][13] ) );
  DFF_X1 \xmem_inst/mem_reg[31][12]  ( .D(n5148), .CK(clk), .QN(
        \xmem_inst/mem[31][12] ) );
  DFF_X1 \xmem_inst/mem_reg[31][10]  ( .D(n5146), .CK(clk), .QN(
        \xmem_inst/mem[31][10] ) );
  DFF_X1 \xmem_inst/mem_reg[31][4]  ( .D(n5140), .CK(clk), .QN(
        \xmem_inst/mem[31][4] ) );
  DFF_X1 \xmem_inst/mem_reg[31][3]  ( .D(n5139), .CK(clk), .QN(
        \xmem_inst/mem[31][3] ) );
  DFF_X1 \xmem_inst/mem_reg[31][2]  ( .D(n5138), .CK(clk), .QN(
        \xmem_inst/mem[31][2] ) );
  DFF_X1 \xmem_inst/mem_reg[31][1]  ( .D(n5137), .CK(clk), .QN(
        \xmem_inst/mem[31][1] ) );
  DFF_X1 \xmem_inst/mem_reg[31][0]  ( .D(n5136), .CK(clk), .QN(
        \xmem_inst/mem[31][0] ) );
  DFF_X1 \xmem_inst/mem_reg[15][28]  ( .D(n4652), .CK(clk), .QN(
        \xmem_inst/mem[15][28] ) );
  DFF_X1 \xmem_inst/mem_reg[15][26]  ( .D(n4650), .CK(clk), .QN(
        \xmem_inst/mem[15][26] ) );
  DFF_X1 \xmem_inst/mem_reg[15][24]  ( .D(n4648), .CK(clk), .QN(
        \xmem_inst/mem[15][24] ) );
  DFF_X1 \xmem_inst/mem_reg[15][23]  ( .D(n4647), .CK(clk), .QN(
        \xmem_inst/mem[15][23] ) );
  DFF_X1 \xmem_inst/mem_reg[15][22]  ( .D(n4646), .CK(clk), .QN(
        \xmem_inst/mem[15][22] ) );
  DFF_X1 \xmem_inst/mem_reg[15][21]  ( .D(n4645), .CK(clk), .QN(
        \xmem_inst/mem[15][21] ) );
  DFF_X1 \xmem_inst/mem_reg[15][20]  ( .D(n4644), .CK(clk), .QN(
        \xmem_inst/mem[15][20] ) );
  DFF_X1 \xmem_inst/mem_reg[15][18]  ( .D(n4642), .CK(clk), .QN(
        \xmem_inst/mem[15][18] ) );
  DFF_X1 \xmem_inst/mem_reg[15][17]  ( .D(n4641), .CK(clk), .QN(
        \xmem_inst/mem[15][17] ) );
  DFF_X1 \xmem_inst/mem_reg[15][16]  ( .D(n4640), .CK(clk), .QN(
        \xmem_inst/mem[15][16] ) );
  DFF_X1 \xmem_inst/mem_reg[15][13]  ( .D(n4637), .CK(clk), .QN(
        \xmem_inst/mem[15][13] ) );
  DFF_X1 \xmem_inst/mem_reg[15][12]  ( .D(n4636), .CK(clk), .QN(
        \xmem_inst/mem[15][12] ) );
  DFF_X1 \xmem_inst/mem_reg[15][10]  ( .D(n4634), .CK(clk), .QN(
        \xmem_inst/mem[15][10] ) );
  DFF_X1 \xmem_inst/mem_reg[15][4]  ( .D(n4628), .CK(clk), .QN(
        \xmem_inst/mem[15][4] ) );
  DFF_X1 \xmem_inst/mem_reg[15][3]  ( .D(n4627), .CK(clk), .QN(
        \xmem_inst/mem[15][3] ) );
  DFF_X1 \xmem_inst/mem_reg[15][2]  ( .D(n4626), .CK(clk), .QN(
        \xmem_inst/mem[15][2] ) );
  DFF_X1 \xmem_inst/mem_reg[15][1]  ( .D(n4625), .CK(clk), .QN(
        \xmem_inst/mem[15][1] ) );
  DFF_X1 \xmem_inst/mem_reg[15][0]  ( .D(n4624), .CK(clk), .QN(
        \xmem_inst/mem[15][0] ) );
  DFF_X1 \xmem_inst/mem_reg[27][28]  ( .D(n5036), .CK(clk), .QN(
        \xmem_inst/mem[27][28] ) );
  DFF_X1 \xmem_inst/mem_reg[27][26]  ( .D(n5034), .CK(clk), .QN(
        \xmem_inst/mem[27][26] ) );
  DFF_X1 \xmem_inst/mem_reg[27][24]  ( .D(n5032), .CK(clk), .QN(
        \xmem_inst/mem[27][24] ) );
  DFF_X1 \xmem_inst/mem_reg[27][23]  ( .D(n5031), .CK(clk), .QN(
        \xmem_inst/mem[27][23] ) );
  DFF_X1 \xmem_inst/mem_reg[27][22]  ( .D(n5030), .CK(clk), .QN(
        \xmem_inst/mem[27][22] ) );
  DFF_X1 \xmem_inst/mem_reg[27][21]  ( .D(n5029), .CK(clk), .QN(
        \xmem_inst/mem[27][21] ) );
  DFF_X1 \xmem_inst/mem_reg[27][20]  ( .D(n5028), .CK(clk), .QN(
        \xmem_inst/mem[27][20] ) );
  DFF_X1 \xmem_inst/mem_reg[27][18]  ( .D(n5026), .CK(clk), .QN(
        \xmem_inst/mem[27][18] ) );
  DFF_X1 \xmem_inst/mem_reg[27][17]  ( .D(n5025), .CK(clk), .QN(
        \xmem_inst/mem[27][17] ) );
  DFF_X1 \xmem_inst/mem_reg[27][16]  ( .D(n5024), .CK(clk), .QN(
        \xmem_inst/mem[27][16] ) );
  DFF_X1 \xmem_inst/mem_reg[27][13]  ( .D(n5021), .CK(clk), .QN(
        \xmem_inst/mem[27][13] ) );
  DFF_X1 \xmem_inst/mem_reg[27][12]  ( .D(n5020), .CK(clk), .QN(
        \xmem_inst/mem[27][12] ) );
  DFF_X1 \xmem_inst/mem_reg[27][10]  ( .D(n5018), .CK(clk), .QN(
        \xmem_inst/mem[27][10] ) );
  DFF_X1 \xmem_inst/mem_reg[27][4]  ( .D(n5012), .CK(clk), .QN(
        \xmem_inst/mem[27][4] ) );
  DFF_X1 \xmem_inst/mem_reg[27][3]  ( .D(n5011), .CK(clk), .QN(
        \xmem_inst/mem[27][3] ) );
  DFF_X1 \xmem_inst/mem_reg[27][2]  ( .D(n5010), .CK(clk), .QN(
        \xmem_inst/mem[27][2] ) );
  DFF_X1 \xmem_inst/mem_reg[27][1]  ( .D(n5009), .CK(clk), .QN(
        \xmem_inst/mem[27][1] ) );
  DFF_X1 \xmem_inst/mem_reg[27][0]  ( .D(n5008), .CK(clk), .QN(
        \xmem_inst/mem[27][0] ) );
  DFF_X1 \xmem_inst/mem_reg[11][28]  ( .D(n4524), .CK(clk), .QN(
        \xmem_inst/mem[11][28] ) );
  DFF_X1 \xmem_inst/mem_reg[11][26]  ( .D(n4522), .CK(clk), .QN(
        \xmem_inst/mem[11][26] ) );
  DFF_X1 \xmem_inst/mem_reg[11][24]  ( .D(n4520), .CK(clk), .QN(
        \xmem_inst/mem[11][24] ) );
  DFF_X1 \xmem_inst/mem_reg[11][23]  ( .D(n4519), .CK(clk), .QN(
        \xmem_inst/mem[11][23] ) );
  DFF_X1 \xmem_inst/mem_reg[11][22]  ( .D(n4518), .CK(clk), .QN(
        \xmem_inst/mem[11][22] ) );
  DFF_X1 \xmem_inst/mem_reg[11][21]  ( .D(n4517), .CK(clk), .QN(
        \xmem_inst/mem[11][21] ) );
  DFF_X1 \xmem_inst/mem_reg[11][20]  ( .D(n4516), .CK(clk), .QN(
        \xmem_inst/mem[11][20] ) );
  DFF_X1 \xmem_inst/mem_reg[11][18]  ( .D(n4514), .CK(clk), .QN(
        \xmem_inst/mem[11][18] ) );
  DFF_X1 \xmem_inst/mem_reg[11][17]  ( .D(n4513), .CK(clk), .QN(
        \xmem_inst/mem[11][17] ) );
  DFF_X1 \xmem_inst/mem_reg[11][16]  ( .D(n4512), .CK(clk), .QN(
        \xmem_inst/mem[11][16] ) );
  DFF_X1 \xmem_inst/mem_reg[11][13]  ( .D(n4509), .CK(clk), .QN(
        \xmem_inst/mem[11][13] ) );
  DFF_X1 \xmem_inst/mem_reg[11][12]  ( .D(n4508), .CK(clk), .QN(
        \xmem_inst/mem[11][12] ) );
  DFF_X1 \xmem_inst/mem_reg[11][10]  ( .D(n4506), .CK(clk), .QN(
        \xmem_inst/mem[11][10] ) );
  DFF_X1 \xmem_inst/mem_reg[11][4]  ( .D(n4500), .CK(clk), .QN(
        \xmem_inst/mem[11][4] ) );
  DFF_X1 \xmem_inst/mem_reg[11][3]  ( .D(n4499), .CK(clk), .QN(
        \xmem_inst/mem[11][3] ) );
  DFF_X1 \xmem_inst/mem_reg[11][2]  ( .D(n4498), .CK(clk), .QN(
        \xmem_inst/mem[11][2] ) );
  DFF_X1 \xmem_inst/mem_reg[11][1]  ( .D(n4497), .CK(clk), .QN(
        \xmem_inst/mem[11][1] ) );
  DFF_X1 \xmem_inst/mem_reg[11][0]  ( .D(n4496), .CK(clk), .QN(
        \xmem_inst/mem[11][0] ) );
  DFF_X1 \xmem_inst/mem_reg[30][28]  ( .D(n5132), .CK(clk), .QN(
        \xmem_inst/mem[30][28] ) );
  DFF_X1 \xmem_inst/mem_reg[30][26]  ( .D(n5130), .CK(clk), .QN(
        \xmem_inst/mem[30][26] ) );
  DFF_X1 \xmem_inst/mem_reg[30][24]  ( .D(n5128), .CK(clk), .QN(
        \xmem_inst/mem[30][24] ) );
  DFF_X1 \xmem_inst/mem_reg[30][23]  ( .D(n5127), .CK(clk), .QN(
        \xmem_inst/mem[30][23] ) );
  DFF_X1 \xmem_inst/mem_reg[30][22]  ( .D(n5126), .CK(clk), .QN(
        \xmem_inst/mem[30][22] ) );
  DFF_X1 \xmem_inst/mem_reg[30][21]  ( .D(n5125), .CK(clk), .QN(
        \xmem_inst/mem[30][21] ) );
  DFF_X1 \xmem_inst/mem_reg[30][20]  ( .D(n5124), .CK(clk), .QN(
        \xmem_inst/mem[30][20] ) );
  DFF_X1 \xmem_inst/mem_reg[30][18]  ( .D(n5122), .CK(clk), .QN(
        \xmem_inst/mem[30][18] ) );
  DFF_X1 \xmem_inst/mem_reg[30][17]  ( .D(n5121), .CK(clk), .QN(
        \xmem_inst/mem[30][17] ) );
  DFF_X1 \xmem_inst/mem_reg[30][16]  ( .D(n5120), .CK(clk), .QN(
        \xmem_inst/mem[30][16] ) );
  DFF_X1 \xmem_inst/mem_reg[30][13]  ( .D(n5117), .CK(clk), .QN(
        \xmem_inst/mem[30][13] ) );
  DFF_X1 \xmem_inst/mem_reg[30][12]  ( .D(n5116), .CK(clk), .QN(
        \xmem_inst/mem[30][12] ) );
  DFF_X1 \xmem_inst/mem_reg[30][10]  ( .D(n5114), .CK(clk), .QN(
        \xmem_inst/mem[30][10] ) );
  DFF_X1 \xmem_inst/mem_reg[30][4]  ( .D(n5108), .CK(clk), .QN(
        \xmem_inst/mem[30][4] ) );
  DFF_X1 \xmem_inst/mem_reg[30][3]  ( .D(n5107), .CK(clk), .QN(
        \xmem_inst/mem[30][3] ) );
  DFF_X1 \xmem_inst/mem_reg[30][2]  ( .D(n5106), .CK(clk), .QN(
        \xmem_inst/mem[30][2] ) );
  DFF_X1 \xmem_inst/mem_reg[30][1]  ( .D(n5105), .CK(clk), .QN(
        \xmem_inst/mem[30][1] ) );
  DFF_X1 \xmem_inst/mem_reg[30][0]  ( .D(n5104), .CK(clk), .QN(
        \xmem_inst/mem[30][0] ) );
  DFF_X1 \xmem_inst/mem_reg[29][28]  ( .D(n5100), .CK(clk), .QN(
        \xmem_inst/mem[29][28] ) );
  DFF_X1 \xmem_inst/mem_reg[29][26]  ( .D(n5098), .CK(clk), .QN(
        \xmem_inst/mem[29][26] ) );
  DFF_X1 \xmem_inst/mem_reg[29][24]  ( .D(n5096), .CK(clk), .QN(
        \xmem_inst/mem[29][24] ) );
  DFF_X1 \xmem_inst/mem_reg[29][23]  ( .D(n5095), .CK(clk), .QN(
        \xmem_inst/mem[29][23] ) );
  DFF_X1 \xmem_inst/mem_reg[29][22]  ( .D(n5094), .CK(clk), .QN(
        \xmem_inst/mem[29][22] ) );
  DFF_X1 \xmem_inst/mem_reg[29][21]  ( .D(n5093), .CK(clk), .QN(
        \xmem_inst/mem[29][21] ) );
  DFF_X1 \xmem_inst/mem_reg[29][20]  ( .D(n5092), .CK(clk), .QN(
        \xmem_inst/mem[29][20] ) );
  DFF_X1 \xmem_inst/mem_reg[29][18]  ( .D(n5090), .CK(clk), .QN(
        \xmem_inst/mem[29][18] ) );
  DFF_X1 \xmem_inst/mem_reg[29][17]  ( .D(n5089), .CK(clk), .QN(
        \xmem_inst/mem[29][17] ) );
  DFF_X1 \xmem_inst/mem_reg[29][16]  ( .D(n5088), .CK(clk), .QN(
        \xmem_inst/mem[29][16] ) );
  DFF_X1 \xmem_inst/mem_reg[29][13]  ( .D(n5085), .CK(clk), .QN(
        \xmem_inst/mem[29][13] ) );
  DFF_X1 \xmem_inst/mem_reg[29][12]  ( .D(n5084), .CK(clk), .QN(
        \xmem_inst/mem[29][12] ) );
  DFF_X1 \xmem_inst/mem_reg[29][10]  ( .D(n5082), .CK(clk), .QN(
        \xmem_inst/mem[29][10] ) );
  DFF_X1 \xmem_inst/mem_reg[29][4]  ( .D(n5076), .CK(clk), .QN(
        \xmem_inst/mem[29][4] ) );
  DFF_X1 \xmem_inst/mem_reg[29][3]  ( .D(n5075), .CK(clk), .QN(
        \xmem_inst/mem[29][3] ) );
  DFF_X1 \xmem_inst/mem_reg[29][2]  ( .D(n5074), .CK(clk), .QN(
        \xmem_inst/mem[29][2] ) );
  DFF_X1 \xmem_inst/mem_reg[29][1]  ( .D(n5073), .CK(clk), .QN(
        \xmem_inst/mem[29][1] ) );
  DFF_X1 \xmem_inst/mem_reg[29][0]  ( .D(n5072), .CK(clk), .QN(
        \xmem_inst/mem[29][0] ) );
  DFF_X1 \xmem_inst/mem_reg[28][28]  ( .D(n5068), .CK(clk), .QN(
        \xmem_inst/mem[28][28] ) );
  DFF_X1 \xmem_inst/mem_reg[28][26]  ( .D(n5066), .CK(clk), .QN(
        \xmem_inst/mem[28][26] ) );
  DFF_X1 \xmem_inst/mem_reg[28][24]  ( .D(n5064), .CK(clk), .QN(
        \xmem_inst/mem[28][24] ) );
  DFF_X1 \xmem_inst/mem_reg[28][23]  ( .D(n5063), .CK(clk), .QN(
        \xmem_inst/mem[28][23] ) );
  DFF_X1 \xmem_inst/mem_reg[28][22]  ( .D(n5062), .CK(clk), .QN(
        \xmem_inst/mem[28][22] ) );
  DFF_X1 \xmem_inst/mem_reg[28][21]  ( .D(n5061), .CK(clk), .QN(
        \xmem_inst/mem[28][21] ) );
  DFF_X1 \xmem_inst/mem_reg[28][20]  ( .D(n5060), .CK(clk), .QN(
        \xmem_inst/mem[28][20] ) );
  DFF_X1 \xmem_inst/mem_reg[28][18]  ( .D(n5058), .CK(clk), .QN(
        \xmem_inst/mem[28][18] ) );
  DFF_X1 \xmem_inst/mem_reg[28][17]  ( .D(n5057), .CK(clk), .QN(
        \xmem_inst/mem[28][17] ) );
  DFF_X1 \xmem_inst/mem_reg[28][16]  ( .D(n5056), .CK(clk), .QN(
        \xmem_inst/mem[28][16] ) );
  DFF_X1 \xmem_inst/mem_reg[28][13]  ( .D(n5053), .CK(clk), .QN(
        \xmem_inst/mem[28][13] ) );
  DFF_X1 \xmem_inst/mem_reg[28][12]  ( .D(n5052), .CK(clk), .QN(
        \xmem_inst/mem[28][12] ) );
  DFF_X1 \xmem_inst/mem_reg[28][10]  ( .D(n5050), .CK(clk), .QN(
        \xmem_inst/mem[28][10] ) );
  DFF_X1 \xmem_inst/mem_reg[28][4]  ( .D(n5044), .CK(clk), .QN(
        \xmem_inst/mem[28][4] ) );
  DFF_X1 \xmem_inst/mem_reg[28][3]  ( .D(n5043), .CK(clk), .QN(
        \xmem_inst/mem[28][3] ) );
  DFF_X1 \xmem_inst/mem_reg[28][2]  ( .D(n5042), .CK(clk), .QN(
        \xmem_inst/mem[28][2] ) );
  DFF_X1 \xmem_inst/mem_reg[28][1]  ( .D(n5041), .CK(clk), .QN(
        \xmem_inst/mem[28][1] ) );
  DFF_X1 \xmem_inst/mem_reg[28][0]  ( .D(n5040), .CK(clk), .QN(
        \xmem_inst/mem[28][0] ) );
  DFF_X1 \xmem_inst/mem_reg[14][28]  ( .D(n4620), .CK(clk), .QN(
        \xmem_inst/mem[14][28] ) );
  DFF_X1 \xmem_inst/mem_reg[14][26]  ( .D(n4618), .CK(clk), .QN(
        \xmem_inst/mem[14][26] ) );
  DFF_X1 \xmem_inst/mem_reg[14][24]  ( .D(n4616), .CK(clk), .QN(
        \xmem_inst/mem[14][24] ) );
  DFF_X1 \xmem_inst/mem_reg[14][23]  ( .D(n4615), .CK(clk), .QN(
        \xmem_inst/mem[14][23] ) );
  DFF_X1 \xmem_inst/mem_reg[14][22]  ( .D(n4614), .CK(clk), .QN(
        \xmem_inst/mem[14][22] ) );
  DFF_X1 \xmem_inst/mem_reg[14][21]  ( .D(n4613), .CK(clk), .QN(
        \xmem_inst/mem[14][21] ) );
  DFF_X1 \xmem_inst/mem_reg[14][20]  ( .D(n4612), .CK(clk), .QN(
        \xmem_inst/mem[14][20] ) );
  DFF_X1 \xmem_inst/mem_reg[14][18]  ( .D(n4610), .CK(clk), .QN(
        \xmem_inst/mem[14][18] ) );
  DFF_X1 \xmem_inst/mem_reg[14][17]  ( .D(n4609), .CK(clk), .QN(
        \xmem_inst/mem[14][17] ) );
  DFF_X1 \xmem_inst/mem_reg[14][16]  ( .D(n4608), .CK(clk), .QN(
        \xmem_inst/mem[14][16] ) );
  DFF_X1 \xmem_inst/mem_reg[14][13]  ( .D(n4605), .CK(clk), .QN(
        \xmem_inst/mem[14][13] ) );
  DFF_X1 \xmem_inst/mem_reg[14][12]  ( .D(n4604), .CK(clk), .QN(
        \xmem_inst/mem[14][12] ) );
  DFF_X1 \xmem_inst/mem_reg[14][10]  ( .D(n4602), .CK(clk), .QN(
        \xmem_inst/mem[14][10] ) );
  DFF_X1 \xmem_inst/mem_reg[14][4]  ( .D(n4596), .CK(clk), .QN(
        \xmem_inst/mem[14][4] ) );
  DFF_X1 \xmem_inst/mem_reg[14][3]  ( .D(n4595), .CK(clk), .QN(
        \xmem_inst/mem[14][3] ) );
  DFF_X1 \xmem_inst/mem_reg[14][2]  ( .D(n4594), .CK(clk), .QN(
        \xmem_inst/mem[14][2] ) );
  DFF_X1 \xmem_inst/mem_reg[14][1]  ( .D(n4593), .CK(clk), .QN(
        \xmem_inst/mem[14][1] ) );
  DFF_X1 \xmem_inst/mem_reg[14][0]  ( .D(n4592), .CK(clk), .QN(
        \xmem_inst/mem[14][0] ) );
  DFF_X1 \xmem_inst/mem_reg[13][28]  ( .D(n4588), .CK(clk), .QN(
        \xmem_inst/mem[13][28] ) );
  DFF_X1 \xmem_inst/mem_reg[13][26]  ( .D(n4586), .CK(clk), .QN(
        \xmem_inst/mem[13][26] ) );
  DFF_X1 \xmem_inst/mem_reg[13][24]  ( .D(n4584), .CK(clk), .QN(
        \xmem_inst/mem[13][24] ) );
  DFF_X1 \xmem_inst/mem_reg[13][23]  ( .D(n4583), .CK(clk), .QN(
        \xmem_inst/mem[13][23] ) );
  DFF_X1 \xmem_inst/mem_reg[13][22]  ( .D(n4582), .CK(clk), .QN(
        \xmem_inst/mem[13][22] ) );
  DFF_X1 \xmem_inst/mem_reg[13][21]  ( .D(n4581), .CK(clk), .QN(
        \xmem_inst/mem[13][21] ) );
  DFF_X1 \xmem_inst/mem_reg[13][20]  ( .D(n4580), .CK(clk), .QN(
        \xmem_inst/mem[13][20] ) );
  DFF_X1 \xmem_inst/mem_reg[13][18]  ( .D(n4578), .CK(clk), .QN(
        \xmem_inst/mem[13][18] ) );
  DFF_X1 \xmem_inst/mem_reg[13][17]  ( .D(n4577), .CK(clk), .QN(
        \xmem_inst/mem[13][17] ) );
  DFF_X1 \xmem_inst/mem_reg[13][16]  ( .D(n4576), .CK(clk), .QN(
        \xmem_inst/mem[13][16] ) );
  DFF_X1 \xmem_inst/mem_reg[13][13]  ( .D(n4573), .CK(clk), .QN(
        \xmem_inst/mem[13][13] ) );
  DFF_X1 \xmem_inst/mem_reg[13][12]  ( .D(n4572), .CK(clk), .QN(
        \xmem_inst/mem[13][12] ) );
  DFF_X1 \xmem_inst/mem_reg[13][10]  ( .D(n4570), .CK(clk), .QN(
        \xmem_inst/mem[13][10] ) );
  DFF_X1 \xmem_inst/mem_reg[13][4]  ( .D(n4564), .CK(clk), .QN(
        \xmem_inst/mem[13][4] ) );
  DFF_X1 \xmem_inst/mem_reg[13][3]  ( .D(n4563), .CK(clk), .QN(
        \xmem_inst/mem[13][3] ) );
  DFF_X1 \xmem_inst/mem_reg[13][2]  ( .D(n4562), .CK(clk), .QN(
        \xmem_inst/mem[13][2] ) );
  DFF_X1 \xmem_inst/mem_reg[13][1]  ( .D(n4561), .CK(clk), .QN(
        \xmem_inst/mem[13][1] ) );
  DFF_X1 \xmem_inst/mem_reg[13][0]  ( .D(n4560), .CK(clk), .QN(
        \xmem_inst/mem[13][0] ) );
  DFF_X1 \xmem_inst/mem_reg[12][28]  ( .D(n4556), .CK(clk), .QN(
        \xmem_inst/mem[12][28] ) );
  DFF_X1 \xmem_inst/mem_reg[12][26]  ( .D(n4554), .CK(clk), .QN(
        \xmem_inst/mem[12][26] ) );
  DFF_X1 \xmem_inst/mem_reg[12][24]  ( .D(n4552), .CK(clk), .QN(
        \xmem_inst/mem[12][24] ) );
  DFF_X1 \xmem_inst/mem_reg[12][23]  ( .D(n4551), .CK(clk), .QN(
        \xmem_inst/mem[12][23] ) );
  DFF_X1 \xmem_inst/mem_reg[12][22]  ( .D(n4550), .CK(clk), .QN(
        \xmem_inst/mem[12][22] ) );
  DFF_X1 \xmem_inst/mem_reg[12][21]  ( .D(n4549), .CK(clk), .QN(
        \xmem_inst/mem[12][21] ) );
  DFF_X1 \xmem_inst/mem_reg[12][20]  ( .D(n4548), .CK(clk), .QN(
        \xmem_inst/mem[12][20] ) );
  DFF_X1 \xmem_inst/mem_reg[12][18]  ( .D(n4546), .CK(clk), .QN(
        \xmem_inst/mem[12][18] ) );
  DFF_X1 \xmem_inst/mem_reg[12][17]  ( .D(n4545), .CK(clk), .QN(
        \xmem_inst/mem[12][17] ) );
  DFF_X1 \xmem_inst/mem_reg[12][16]  ( .D(n4544), .CK(clk), .QN(
        \xmem_inst/mem[12][16] ) );
  DFF_X1 \xmem_inst/mem_reg[12][13]  ( .D(n4541), .CK(clk), .QN(
        \xmem_inst/mem[12][13] ) );
  DFF_X1 \xmem_inst/mem_reg[12][12]  ( .D(n4540), .CK(clk), .QN(
        \xmem_inst/mem[12][12] ) );
  DFF_X1 \xmem_inst/mem_reg[12][10]  ( .D(n4538), .CK(clk), .QN(
        \xmem_inst/mem[12][10] ) );
  DFF_X1 \xmem_inst/mem_reg[12][4]  ( .D(n4532), .CK(clk), .QN(
        \xmem_inst/mem[12][4] ) );
  DFF_X1 \xmem_inst/mem_reg[12][3]  ( .D(n4531), .CK(clk), .QN(
        \xmem_inst/mem[12][3] ) );
  DFF_X1 \xmem_inst/mem_reg[12][2]  ( .D(n4530), .CK(clk), .QN(
        \xmem_inst/mem[12][2] ) );
  DFF_X1 \xmem_inst/mem_reg[12][1]  ( .D(n4529), .CK(clk), .QN(
        \xmem_inst/mem[12][1] ) );
  DFF_X1 \xmem_inst/mem_reg[12][0]  ( .D(n4528), .CK(clk), .QN(
        \xmem_inst/mem[12][0] ) );
  DFF_X1 \xmem_inst/mem_reg[26][28]  ( .D(n5004), .CK(clk), .QN(
        \xmem_inst/mem[26][28] ) );
  DFF_X1 \xmem_inst/mem_reg[26][26]  ( .D(n5002), .CK(clk), .QN(
        \xmem_inst/mem[26][26] ) );
  DFF_X1 \xmem_inst/mem_reg[26][24]  ( .D(n5000), .CK(clk), .QN(
        \xmem_inst/mem[26][24] ) );
  DFF_X1 \xmem_inst/mem_reg[26][23]  ( .D(n4999), .CK(clk), .QN(
        \xmem_inst/mem[26][23] ) );
  DFF_X1 \xmem_inst/mem_reg[26][22]  ( .D(n4998), .CK(clk), .QN(
        \xmem_inst/mem[26][22] ) );
  DFF_X1 \xmem_inst/mem_reg[26][21]  ( .D(n4997), .CK(clk), .QN(
        \xmem_inst/mem[26][21] ) );
  DFF_X1 \xmem_inst/mem_reg[26][20]  ( .D(n4996), .CK(clk), .QN(
        \xmem_inst/mem[26][20] ) );
  DFF_X1 \xmem_inst/mem_reg[26][18]  ( .D(n4994), .CK(clk), .QN(
        \xmem_inst/mem[26][18] ) );
  DFF_X1 \xmem_inst/mem_reg[26][17]  ( .D(n4993), .CK(clk), .QN(
        \xmem_inst/mem[26][17] ) );
  DFF_X1 \xmem_inst/mem_reg[26][16]  ( .D(n4992), .CK(clk), .QN(
        \xmem_inst/mem[26][16] ) );
  DFF_X1 \xmem_inst/mem_reg[26][13]  ( .D(n4989), .CK(clk), .QN(
        \xmem_inst/mem[26][13] ) );
  DFF_X1 \xmem_inst/mem_reg[26][12]  ( .D(n4988), .CK(clk), .QN(
        \xmem_inst/mem[26][12] ) );
  DFF_X1 \xmem_inst/mem_reg[26][10]  ( .D(n4986), .CK(clk), .QN(
        \xmem_inst/mem[26][10] ) );
  DFF_X1 \xmem_inst/mem_reg[26][4]  ( .D(n4980), .CK(clk), .QN(
        \xmem_inst/mem[26][4] ) );
  DFF_X1 \xmem_inst/mem_reg[26][3]  ( .D(n4979), .CK(clk), .QN(
        \xmem_inst/mem[26][3] ) );
  DFF_X1 \xmem_inst/mem_reg[26][2]  ( .D(n4978), .CK(clk), .QN(
        \xmem_inst/mem[26][2] ) );
  DFF_X1 \xmem_inst/mem_reg[26][1]  ( .D(n4977), .CK(clk), .QN(
        \xmem_inst/mem[26][1] ) );
  DFF_X1 \xmem_inst/mem_reg[26][0]  ( .D(n4976), .CK(clk), .QN(
        \xmem_inst/mem[26][0] ) );
  DFF_X1 \xmem_inst/mem_reg[10][28]  ( .D(n4492), .CK(clk), .QN(
        \xmem_inst/mem[10][28] ) );
  DFF_X1 \xmem_inst/mem_reg[10][26]  ( .D(n4490), .CK(clk), .QN(
        \xmem_inst/mem[10][26] ) );
  DFF_X1 \xmem_inst/mem_reg[10][24]  ( .D(n4488), .CK(clk), .QN(
        \xmem_inst/mem[10][24] ) );
  DFF_X1 \xmem_inst/mem_reg[10][23]  ( .D(n4487), .CK(clk), .QN(
        \xmem_inst/mem[10][23] ) );
  DFF_X1 \xmem_inst/mem_reg[10][22]  ( .D(n4486), .CK(clk), .QN(
        \xmem_inst/mem[10][22] ) );
  DFF_X1 \xmem_inst/mem_reg[10][21]  ( .D(n4485), .CK(clk), .QN(
        \xmem_inst/mem[10][21] ) );
  DFF_X1 \xmem_inst/mem_reg[10][20]  ( .D(n4484), .CK(clk), .QN(
        \xmem_inst/mem[10][20] ) );
  DFF_X1 \xmem_inst/mem_reg[10][18]  ( .D(n4482), .CK(clk), .QN(
        \xmem_inst/mem[10][18] ) );
  DFF_X1 \xmem_inst/mem_reg[10][17]  ( .D(n4481), .CK(clk), .QN(
        \xmem_inst/mem[10][17] ) );
  DFF_X1 \xmem_inst/mem_reg[10][16]  ( .D(n4480), .CK(clk), .QN(
        \xmem_inst/mem[10][16] ) );
  DFF_X1 \xmem_inst/mem_reg[10][13]  ( .D(n4477), .CK(clk), .QN(
        \xmem_inst/mem[10][13] ) );
  DFF_X1 \xmem_inst/mem_reg[10][12]  ( .D(n4476), .CK(clk), .QN(
        \xmem_inst/mem[10][12] ) );
  DFF_X1 \xmem_inst/mem_reg[10][10]  ( .D(n4474), .CK(clk), .QN(
        \xmem_inst/mem[10][10] ) );
  DFF_X1 \xmem_inst/mem_reg[10][4]  ( .D(n4468), .CK(clk), .QN(
        \xmem_inst/mem[10][4] ) );
  DFF_X1 \xmem_inst/mem_reg[10][3]  ( .D(n4467), .CK(clk), .QN(
        \xmem_inst/mem[10][3] ) );
  DFF_X1 \xmem_inst/mem_reg[10][2]  ( .D(n4466), .CK(clk), .QN(
        \xmem_inst/mem[10][2] ) );
  DFF_X1 \xmem_inst/mem_reg[10][1]  ( .D(n4465), .CK(clk), .QN(
        \xmem_inst/mem[10][1] ) );
  DFF_X1 \xmem_inst/mem_reg[10][0]  ( .D(n4464), .CK(clk), .QN(
        \xmem_inst/mem[10][0] ) );
  DFF_X1 \xmem_inst/mem_reg[25][28]  ( .D(n4972), .CK(clk), .QN(
        \xmem_inst/mem[25][28] ) );
  DFF_X1 \xmem_inst/mem_reg[25][26]  ( .D(n4970), .CK(clk), .QN(
        \xmem_inst/mem[25][26] ) );
  DFF_X1 \xmem_inst/mem_reg[25][24]  ( .D(n4968), .CK(clk), .QN(
        \xmem_inst/mem[25][24] ) );
  DFF_X1 \xmem_inst/mem_reg[25][23]  ( .D(n4967), .CK(clk), .QN(
        \xmem_inst/mem[25][23] ) );
  DFF_X1 \xmem_inst/mem_reg[25][22]  ( .D(n4966), .CK(clk), .QN(
        \xmem_inst/mem[25][22] ) );
  DFF_X1 \xmem_inst/mem_reg[25][21]  ( .D(n4965), .CK(clk), .QN(
        \xmem_inst/mem[25][21] ) );
  DFF_X1 \xmem_inst/mem_reg[25][20]  ( .D(n4964), .CK(clk), .QN(
        \xmem_inst/mem[25][20] ) );
  DFF_X1 \xmem_inst/mem_reg[25][18]  ( .D(n4962), .CK(clk), .QN(
        \xmem_inst/mem[25][18] ) );
  DFF_X1 \xmem_inst/mem_reg[25][17]  ( .D(n4961), .CK(clk), .QN(
        \xmem_inst/mem[25][17] ) );
  DFF_X1 \xmem_inst/mem_reg[25][16]  ( .D(n4960), .CK(clk), .QN(
        \xmem_inst/mem[25][16] ) );
  DFF_X1 \xmem_inst/mem_reg[25][13]  ( .D(n4957), .CK(clk), .QN(
        \xmem_inst/mem[25][13] ) );
  DFF_X1 \xmem_inst/mem_reg[25][12]  ( .D(n4956), .CK(clk), .QN(
        \xmem_inst/mem[25][12] ) );
  DFF_X1 \xmem_inst/mem_reg[25][10]  ( .D(n4954), .CK(clk), .QN(
        \xmem_inst/mem[25][10] ) );
  DFF_X1 \xmem_inst/mem_reg[25][4]  ( .D(n4948), .CK(clk), .QN(
        \xmem_inst/mem[25][4] ) );
  DFF_X1 \xmem_inst/mem_reg[25][3]  ( .D(n4947), .CK(clk), .QN(
        \xmem_inst/mem[25][3] ) );
  DFF_X1 \xmem_inst/mem_reg[25][2]  ( .D(n4946), .CK(clk), .QN(
        \xmem_inst/mem[25][2] ) );
  DFF_X1 \xmem_inst/mem_reg[25][1]  ( .D(n4945), .CK(clk), .QN(
        \xmem_inst/mem[25][1] ) );
  DFF_X1 \xmem_inst/mem_reg[25][0]  ( .D(n4944), .CK(clk), .QN(
        \xmem_inst/mem[25][0] ) );
  DFF_X1 \xmem_inst/mem_reg[24][28]  ( .D(n4940), .CK(clk), .QN(
        \xmem_inst/mem[24][28] ) );
  DFF_X1 \xmem_inst/mem_reg[24][26]  ( .D(n4938), .CK(clk), .QN(
        \xmem_inst/mem[24][26] ) );
  DFF_X1 \xmem_inst/mem_reg[24][24]  ( .D(n4936), .CK(clk), .QN(
        \xmem_inst/mem[24][24] ) );
  DFF_X1 \xmem_inst/mem_reg[24][23]  ( .D(n4935), .CK(clk), .QN(
        \xmem_inst/mem[24][23] ) );
  DFF_X1 \xmem_inst/mem_reg[24][22]  ( .D(n4934), .CK(clk), .QN(
        \xmem_inst/mem[24][22] ) );
  DFF_X1 \xmem_inst/mem_reg[24][21]  ( .D(n4933), .CK(clk), .QN(
        \xmem_inst/mem[24][21] ) );
  DFF_X1 \xmem_inst/mem_reg[24][20]  ( .D(n4932), .CK(clk), .QN(
        \xmem_inst/mem[24][20] ) );
  DFF_X1 \xmem_inst/mem_reg[24][18]  ( .D(n4930), .CK(clk), .QN(
        \xmem_inst/mem[24][18] ) );
  DFF_X1 \xmem_inst/mem_reg[24][17]  ( .D(n4929), .CK(clk), .QN(
        \xmem_inst/mem[24][17] ) );
  DFF_X1 \xmem_inst/mem_reg[24][16]  ( .D(n4928), .CK(clk), .QN(
        \xmem_inst/mem[24][16] ) );
  DFF_X1 \xmem_inst/mem_reg[24][13]  ( .D(n4925), .CK(clk), .QN(
        \xmem_inst/mem[24][13] ) );
  DFF_X1 \xmem_inst/mem_reg[24][12]  ( .D(n4924), .CK(clk), .QN(
        \xmem_inst/mem[24][12] ) );
  DFF_X1 \xmem_inst/mem_reg[24][10]  ( .D(n4922), .CK(clk), .QN(
        \xmem_inst/mem[24][10] ) );
  DFF_X1 \xmem_inst/mem_reg[24][4]  ( .D(n4916), .CK(clk), .QN(
        \xmem_inst/mem[24][4] ) );
  DFF_X1 \xmem_inst/mem_reg[24][3]  ( .D(n4915), .CK(clk), .QN(
        \xmem_inst/mem[24][3] ) );
  DFF_X1 \xmem_inst/mem_reg[24][2]  ( .D(n4914), .CK(clk), .QN(
        \xmem_inst/mem[24][2] ) );
  DFF_X1 \xmem_inst/mem_reg[24][1]  ( .D(n4913), .CK(clk), .QN(
        \xmem_inst/mem[24][1] ) );
  DFF_X1 \xmem_inst/mem_reg[24][0]  ( .D(n4912), .CK(clk), .QN(
        \xmem_inst/mem[24][0] ) );
  DFF_X1 \xmem_inst/mem_reg[9][28]  ( .D(n4460), .CK(clk), .QN(
        \xmem_inst/mem[9][28] ) );
  DFF_X1 \xmem_inst/mem_reg[9][26]  ( .D(n4458), .CK(clk), .QN(
        \xmem_inst/mem[9][26] ) );
  DFF_X1 \xmem_inst/mem_reg[9][24]  ( .D(n4456), .CK(clk), .QN(
        \xmem_inst/mem[9][24] ) );
  DFF_X1 \xmem_inst/mem_reg[9][23]  ( .D(n4455), .CK(clk), .QN(
        \xmem_inst/mem[9][23] ) );
  DFF_X1 \xmem_inst/mem_reg[9][22]  ( .D(n4454), .CK(clk), .QN(
        \xmem_inst/mem[9][22] ) );
  DFF_X1 \xmem_inst/mem_reg[9][21]  ( .D(n4453), .CK(clk), .QN(
        \xmem_inst/mem[9][21] ) );
  DFF_X1 \xmem_inst/mem_reg[9][20]  ( .D(n4452), .CK(clk), .QN(
        \xmem_inst/mem[9][20] ) );
  DFF_X1 \xmem_inst/mem_reg[9][18]  ( .D(n4450), .CK(clk), .QN(
        \xmem_inst/mem[9][18] ) );
  DFF_X1 \xmem_inst/mem_reg[9][17]  ( .D(n4449), .CK(clk), .QN(
        \xmem_inst/mem[9][17] ) );
  DFF_X1 \xmem_inst/mem_reg[9][16]  ( .D(n4448), .CK(clk), .QN(
        \xmem_inst/mem[9][16] ) );
  DFF_X1 \xmem_inst/mem_reg[9][13]  ( .D(n4445), .CK(clk), .QN(
        \xmem_inst/mem[9][13] ) );
  DFF_X1 \xmem_inst/mem_reg[9][12]  ( .D(n4444), .CK(clk), .QN(
        \xmem_inst/mem[9][12] ) );
  DFF_X1 \xmem_inst/mem_reg[9][10]  ( .D(n4442), .CK(clk), .QN(
        \xmem_inst/mem[9][10] ) );
  DFF_X1 \xmem_inst/mem_reg[9][4]  ( .D(n4436), .CK(clk), .QN(
        \xmem_inst/mem[9][4] ) );
  DFF_X1 \xmem_inst/mem_reg[9][3]  ( .D(n4435), .CK(clk), .QN(
        \xmem_inst/mem[9][3] ) );
  DFF_X1 \xmem_inst/mem_reg[9][2]  ( .D(n4434), .CK(clk), .QN(
        \xmem_inst/mem[9][2] ) );
  DFF_X1 \xmem_inst/mem_reg[9][1]  ( .D(n4433), .CK(clk), .QN(
        \xmem_inst/mem[9][1] ) );
  DFF_X1 \xmem_inst/mem_reg[9][0]  ( .D(n4432), .CK(clk), .QN(
        \xmem_inst/mem[9][0] ) );
  DFF_X1 \xmem_inst/mem_reg[8][28]  ( .D(n4428), .CK(clk), .QN(
        \xmem_inst/mem[8][28] ) );
  DFF_X1 \xmem_inst/mem_reg[8][26]  ( .D(n4426), .CK(clk), .QN(
        \xmem_inst/mem[8][26] ) );
  DFF_X1 \xmem_inst/mem_reg[8][24]  ( .D(n4424), .CK(clk), .QN(
        \xmem_inst/mem[8][24] ) );
  DFF_X1 \xmem_inst/mem_reg[8][23]  ( .D(n4423), .CK(clk), .QN(
        \xmem_inst/mem[8][23] ) );
  DFF_X1 \xmem_inst/mem_reg[8][22]  ( .D(n4422), .CK(clk), .QN(
        \xmem_inst/mem[8][22] ) );
  DFF_X1 \xmem_inst/mem_reg[8][21]  ( .D(n4421), .CK(clk), .QN(
        \xmem_inst/mem[8][21] ) );
  DFF_X1 \xmem_inst/mem_reg[8][20]  ( .D(n4420), .CK(clk), .QN(
        \xmem_inst/mem[8][20] ) );
  DFF_X1 \xmem_inst/mem_reg[8][18]  ( .D(n4418), .CK(clk), .QN(
        \xmem_inst/mem[8][18] ) );
  DFF_X1 \xmem_inst/mem_reg[8][17]  ( .D(n4417), .CK(clk), .QN(
        \xmem_inst/mem[8][17] ) );
  DFF_X1 \xmem_inst/mem_reg[8][16]  ( .D(n4416), .CK(clk), .QN(
        \xmem_inst/mem[8][16] ) );
  DFF_X1 \xmem_inst/mem_reg[8][13]  ( .D(n4413), .CK(clk), .QN(
        \xmem_inst/mem[8][13] ) );
  DFF_X1 \xmem_inst/mem_reg[8][12]  ( .D(n4412), .CK(clk), .QN(
        \xmem_inst/mem[8][12] ) );
  DFF_X1 \xmem_inst/mem_reg[8][10]  ( .D(n4410), .CK(clk), .QN(
        \xmem_inst/mem[8][10] ) );
  DFF_X1 \xmem_inst/mem_reg[8][4]  ( .D(n4404), .CK(clk), .QN(
        \xmem_inst/mem[8][4] ) );
  DFF_X1 \xmem_inst/mem_reg[8][3]  ( .D(n4403), .CK(clk), .QN(
        \xmem_inst/mem[8][3] ) );
  DFF_X1 \xmem_inst/mem_reg[8][2]  ( .D(n4402), .CK(clk), .QN(
        \xmem_inst/mem[8][2] ) );
  DFF_X1 \xmem_inst/mem_reg[8][1]  ( .D(n4401), .CK(clk), .QN(
        \xmem_inst/mem[8][1] ) );
  DFF_X1 \xmem_inst/mem_reg[8][0]  ( .D(n4400), .CK(clk), .QN(
        \xmem_inst/mem[8][0] ) );
  DFF_X1 \xmem_inst/mem_reg[26][29]  ( .D(n5005), .CK(clk), .QN(
        \xmem_inst/mem[26][29] ) );
  DFF_X1 \xmem_inst/mem_reg[26][27]  ( .D(n5003), .CK(clk), .QN(
        \xmem_inst/mem[26][27] ) );
  DFF_X1 \xmem_inst/mem_reg[26][25]  ( .D(n5001), .CK(clk), .QN(
        \xmem_inst/mem[26][25] ) );
  DFF_X1 \xmem_inst/mem_reg[26][14]  ( .D(n4990), .CK(clk), .QN(
        \xmem_inst/mem[26][14] ) );
  DFF_X1 \xmem_inst/mem_reg[26][11]  ( .D(n4987), .CK(clk), .QN(
        \xmem_inst/mem[26][11] ) );
  DFF_X1 \xmem_inst/mem_reg[26][9]  ( .D(n4985), .CK(clk), .QN(
        \xmem_inst/mem[26][9] ) );
  DFF_X1 \xmem_inst/mem_reg[26][8]  ( .D(n4984), .CK(clk), .QN(
        \xmem_inst/mem[26][8] ) );
  DFF_X1 \xmem_inst/mem_reg[26][7]  ( .D(n4983), .CK(clk), .QN(
        \xmem_inst/mem[26][7] ) );
  DFF_X1 \xmem_inst/mem_reg[26][6]  ( .D(n4982), .CK(clk), .QN(
        \xmem_inst/mem[26][6] ) );
  DFF_X1 \xmem_inst/mem_reg[26][5]  ( .D(n4981), .CK(clk), .QN(
        \xmem_inst/mem[26][5] ) );
  DFF_X1 \xmem_inst/mem_reg[10][29]  ( .D(n4493), .CK(clk), .QN(
        \xmem_inst/mem[10][29] ) );
  DFF_X1 \xmem_inst/mem_reg[10][27]  ( .D(n4491), .CK(clk), .QN(
        \xmem_inst/mem[10][27] ) );
  DFF_X1 \xmem_inst/mem_reg[10][25]  ( .D(n4489), .CK(clk), .QN(
        \xmem_inst/mem[10][25] ) );
  DFF_X1 \xmem_inst/mem_reg[10][14]  ( .D(n4478), .CK(clk), .QN(
        \xmem_inst/mem[10][14] ) );
  DFF_X1 \xmem_inst/mem_reg[10][11]  ( .D(n4475), .CK(clk), .QN(
        \xmem_inst/mem[10][11] ) );
  DFF_X1 \xmem_inst/mem_reg[10][9]  ( .D(n4473), .CK(clk), .QN(
        \xmem_inst/mem[10][9] ) );
  DFF_X1 \xmem_inst/mem_reg[10][8]  ( .D(n4472), .CK(clk), .QN(
        \xmem_inst/mem[10][8] ) );
  DFF_X1 \xmem_inst/mem_reg[10][7]  ( .D(n4471), .CK(clk), .QN(
        \xmem_inst/mem[10][7] ) );
  DFF_X1 \xmem_inst/mem_reg[10][6]  ( .D(n4470), .CK(clk), .QN(
        \xmem_inst/mem[10][6] ) );
  DFF_X1 \xmem_inst/mem_reg[10][5]  ( .D(n4469), .CK(clk), .QN(
        \xmem_inst/mem[10][5] ) );
  DFF_X1 \xmem_inst/mem_reg[25][29]  ( .D(n4973), .CK(clk), .QN(
        \xmem_inst/mem[25][29] ) );
  DFF_X1 \xmem_inst/mem_reg[25][27]  ( .D(n4971), .CK(clk), .QN(
        \xmem_inst/mem[25][27] ) );
  DFF_X1 \xmem_inst/mem_reg[25][25]  ( .D(n4969), .CK(clk), .QN(
        \xmem_inst/mem[25][25] ) );
  DFF_X1 \xmem_inst/mem_reg[25][14]  ( .D(n4958), .CK(clk), .QN(
        \xmem_inst/mem[25][14] ) );
  DFF_X1 \xmem_inst/mem_reg[25][11]  ( .D(n4955), .CK(clk), .QN(
        \xmem_inst/mem[25][11] ) );
  DFF_X1 \xmem_inst/mem_reg[25][9]  ( .D(n4953), .CK(clk), .QN(
        \xmem_inst/mem[25][9] ) );
  DFF_X1 \xmem_inst/mem_reg[25][8]  ( .D(n4952), .CK(clk), .QN(
        \xmem_inst/mem[25][8] ) );
  DFF_X1 \xmem_inst/mem_reg[25][7]  ( .D(n4951), .CK(clk), .QN(
        \xmem_inst/mem[25][7] ) );
  DFF_X1 \xmem_inst/mem_reg[25][6]  ( .D(n4950), .CK(clk), .QN(
        \xmem_inst/mem[25][6] ) );
  DFF_X1 \xmem_inst/mem_reg[25][5]  ( .D(n4949), .CK(clk), .QN(
        \xmem_inst/mem[25][5] ) );
  DFF_X1 \xmem_inst/mem_reg[24][29]  ( .D(n4941), .CK(clk), .QN(
        \xmem_inst/mem[24][29] ) );
  DFF_X1 \xmem_inst/mem_reg[24][27]  ( .D(n4939), .CK(clk), .QN(
        \xmem_inst/mem[24][27] ) );
  DFF_X1 \xmem_inst/mem_reg[24][25]  ( .D(n4937), .CK(clk), .QN(
        \xmem_inst/mem[24][25] ) );
  DFF_X1 \xmem_inst/mem_reg[24][14]  ( .D(n4926), .CK(clk), .QN(
        \xmem_inst/mem[24][14] ) );
  DFF_X1 \xmem_inst/mem_reg[24][11]  ( .D(n4923), .CK(clk), .QN(
        \xmem_inst/mem[24][11] ) );
  DFF_X1 \xmem_inst/mem_reg[24][9]  ( .D(n4921), .CK(clk), .QN(
        \xmem_inst/mem[24][9] ) );
  DFF_X1 \xmem_inst/mem_reg[24][8]  ( .D(n4920), .CK(clk), .QN(
        \xmem_inst/mem[24][8] ) );
  DFF_X1 \xmem_inst/mem_reg[24][7]  ( .D(n4919), .CK(clk), .QN(
        \xmem_inst/mem[24][7] ) );
  DFF_X1 \xmem_inst/mem_reg[24][6]  ( .D(n4918), .CK(clk), .QN(
        \xmem_inst/mem[24][6] ) );
  DFF_X1 \xmem_inst/mem_reg[24][5]  ( .D(n4917), .CK(clk), .QN(
        \xmem_inst/mem[24][5] ) );
  DFF_X1 \xmem_inst/mem_reg[9][29]  ( .D(n4461), .CK(clk), .QN(
        \xmem_inst/mem[9][29] ) );
  DFF_X1 \xmem_inst/mem_reg[9][27]  ( .D(n4459), .CK(clk), .QN(
        \xmem_inst/mem[9][27] ) );
  DFF_X1 \xmem_inst/mem_reg[9][25]  ( .D(n4457), .CK(clk), .QN(
        \xmem_inst/mem[9][25] ) );
  DFF_X1 \xmem_inst/mem_reg[9][14]  ( .D(n4446), .CK(clk), .QN(
        \xmem_inst/mem[9][14] ) );
  DFF_X1 \xmem_inst/mem_reg[9][11]  ( .D(n4443), .CK(clk), .QN(
        \xmem_inst/mem[9][11] ) );
  DFF_X1 \xmem_inst/mem_reg[9][9]  ( .D(n4441), .CK(clk), .QN(
        \xmem_inst/mem[9][9] ) );
  DFF_X1 \xmem_inst/mem_reg[9][8]  ( .D(n4440), .CK(clk), .QN(
        \xmem_inst/mem[9][8] ) );
  DFF_X1 \xmem_inst/mem_reg[9][7]  ( .D(n4439), .CK(clk), .QN(
        \xmem_inst/mem[9][7] ) );
  DFF_X1 \xmem_inst/mem_reg[9][6]  ( .D(n4438), .CK(clk), .QN(
        \xmem_inst/mem[9][6] ) );
  DFF_X1 \xmem_inst/mem_reg[9][5]  ( .D(n4437), .CK(clk), .QN(
        \xmem_inst/mem[9][5] ) );
  DFF_X1 \xmem_inst/mem_reg[8][29]  ( .D(n4429), .CK(clk), .QN(
        \xmem_inst/mem[8][29] ) );
  DFF_X1 \xmem_inst/mem_reg[8][27]  ( .D(n4427), .CK(clk), .QN(
        \xmem_inst/mem[8][27] ) );
  DFF_X1 \xmem_inst/mem_reg[8][25]  ( .D(n4425), .CK(clk), .QN(
        \xmem_inst/mem[8][25] ) );
  DFF_X1 \xmem_inst/mem_reg[8][14]  ( .D(n4414), .CK(clk), .QN(
        \xmem_inst/mem[8][14] ) );
  DFF_X1 \xmem_inst/mem_reg[8][11]  ( .D(n4411), .CK(clk), .QN(
        \xmem_inst/mem[8][11] ) );
  DFF_X1 \xmem_inst/mem_reg[8][9]  ( .D(n4409), .CK(clk), .QN(
        \xmem_inst/mem[8][9] ) );
  DFF_X1 \xmem_inst/mem_reg[8][8]  ( .D(n4408), .CK(clk), .QN(
        \xmem_inst/mem[8][8] ) );
  DFF_X1 \xmem_inst/mem_reg[8][7]  ( .D(n4407), .CK(clk), .QN(
        \xmem_inst/mem[8][7] ) );
  DFF_X1 \xmem_inst/mem_reg[8][6]  ( .D(n4406), .CK(clk), .QN(
        \xmem_inst/mem[8][6] ) );
  DFF_X1 \xmem_inst/mem_reg[8][5]  ( .D(n4405), .CK(clk), .QN(
        \xmem_inst/mem[8][5] ) );
  DFF_X1 \xmem_inst/mem_reg[38][31]  ( .D(n5331), .CK(clk), .QN(
        \xmem_inst/mem[38][31] ) );
  DFF_X1 \xmem_inst/mem_reg[38][30]  ( .D(n5330), .CK(clk), .QN(
        \xmem_inst/mem[38][30] ) );
  DFF_X1 \xmem_inst/mem_reg[38][19]  ( .D(n5319), .CK(clk), .QN(
        \xmem_inst/mem[38][19] ) );
  DFF_X1 \xmem_inst/mem_reg[38][16]  ( .D(n5316), .CK(clk), .QN(
        \xmem_inst/mem[38][16] ) );
  DFF_X1 \xmem_inst/mem_reg[37][31]  ( .D(n5299), .CK(clk), .QN(
        \xmem_inst/mem[37][31] ) );
  DFF_X1 \xmem_inst/mem_reg[37][30]  ( .D(n5298), .CK(clk), .QN(
        \xmem_inst/mem[37][30] ) );
  DFF_X1 \xmem_inst/mem_reg[37][19]  ( .D(n5287), .CK(clk), .QN(
        \xmem_inst/mem[37][19] ) );
  DFF_X1 \xmem_inst/mem_reg[37][16]  ( .D(n5284), .CK(clk), .QN(
        \xmem_inst/mem[37][16] ) );
  DFF_X1 \xmem_inst/mem_reg[36][31]  ( .D(n5267), .CK(clk), .QN(
        \xmem_inst/mem[36][31] ) );
  DFF_X1 \xmem_inst/mem_reg[36][30]  ( .D(n5266), .CK(clk), .QN(
        \xmem_inst/mem[36][30] ) );
  DFF_X1 \xmem_inst/mem_reg[36][19]  ( .D(n5255), .CK(clk), .QN(
        \xmem_inst/mem[36][19] ) );
  DFF_X1 \xmem_inst/mem_reg[36][16]  ( .D(n5252), .CK(clk), .QN(
        \xmem_inst/mem[36][16] ) );
  DFF_X1 \xmem_inst/mem_reg[35][31]  ( .D(n5235), .CK(clk), .QN(
        \xmem_inst/mem[35][31] ) );
  DFF_X1 \xmem_inst/mem_reg[35][30]  ( .D(n5234), .CK(clk), .QN(
        \xmem_inst/mem[35][30] ) );
  DFF_X1 \xmem_inst/mem_reg[35][19]  ( .D(n5223), .CK(clk), .QN(
        \xmem_inst/mem[35][19] ) );
  DFF_X1 \xmem_inst/mem_reg[35][16]  ( .D(n5220), .CK(clk), .QN(
        \xmem_inst/mem[35][16] ) );
  DFF_X1 \xmem_inst/mem_reg[38][29]  ( .D(n5329), .CK(clk), .QN(
        \xmem_inst/mem[38][29] ) );
  DFF_X1 \xmem_inst/mem_reg[38][27]  ( .D(n5327), .CK(clk), .QN(
        \xmem_inst/mem[38][27] ) );
  DFF_X1 \xmem_inst/mem_reg[38][25]  ( .D(n5325), .CK(clk), .QN(
        \xmem_inst/mem[38][25] ) );
  DFF_X1 \xmem_inst/mem_reg[38][14]  ( .D(n5314), .CK(clk), .QN(
        \xmem_inst/mem[38][14] ) );
  DFF_X1 \xmem_inst/mem_reg[38][11]  ( .D(n5311), .CK(clk), .QN(
        \xmem_inst/mem[38][11] ) );
  DFF_X1 \xmem_inst/mem_reg[38][9]  ( .D(n5309), .CK(clk), .QN(
        \xmem_inst/mem[38][9] ) );
  DFF_X1 \xmem_inst/mem_reg[38][8]  ( .D(n5308), .CK(clk), .QN(
        \xmem_inst/mem[38][8] ) );
  DFF_X1 \xmem_inst/mem_reg[38][7]  ( .D(n5307), .CK(clk), .QN(
        \xmem_inst/mem[38][7] ) );
  DFF_X1 \xmem_inst/mem_reg[38][6]  ( .D(n5306), .CK(clk), .QN(
        \xmem_inst/mem[38][6] ) );
  DFF_X1 \xmem_inst/mem_reg[38][5]  ( .D(n5305), .CK(clk), .QN(
        \xmem_inst/mem[38][5] ) );
  DFF_X1 \xmem_inst/mem_reg[37][29]  ( .D(n5297), .CK(clk), .QN(
        \xmem_inst/mem[37][29] ) );
  DFF_X1 \xmem_inst/mem_reg[37][27]  ( .D(n5295), .CK(clk), .QN(
        \xmem_inst/mem[37][27] ) );
  DFF_X1 \xmem_inst/mem_reg[37][25]  ( .D(n5293), .CK(clk), .QN(
        \xmem_inst/mem[37][25] ) );
  DFF_X1 \xmem_inst/mem_reg[37][14]  ( .D(n5282), .CK(clk), .QN(
        \xmem_inst/mem[37][14] ) );
  DFF_X1 \xmem_inst/mem_reg[37][11]  ( .D(n5279), .CK(clk), .QN(
        \xmem_inst/mem[37][11] ) );
  DFF_X1 \xmem_inst/mem_reg[37][9]  ( .D(n5277), .CK(clk), .QN(
        \xmem_inst/mem[37][9] ) );
  DFF_X1 \xmem_inst/mem_reg[37][8]  ( .D(n5276), .CK(clk), .QN(
        \xmem_inst/mem[37][8] ) );
  DFF_X1 \xmem_inst/mem_reg[37][7]  ( .D(n5275), .CK(clk), .QN(
        \xmem_inst/mem[37][7] ) );
  DFF_X1 \xmem_inst/mem_reg[37][6]  ( .D(n5274), .CK(clk), .QN(
        \xmem_inst/mem[37][6] ) );
  DFF_X1 \xmem_inst/mem_reg[37][5]  ( .D(n5273), .CK(clk), .QN(
        \xmem_inst/mem[37][5] ) );
  DFF_X1 \xmem_inst/mem_reg[36][29]  ( .D(n5265), .CK(clk), .QN(
        \xmem_inst/mem[36][29] ) );
  DFF_X1 \xmem_inst/mem_reg[36][27]  ( .D(n5263), .CK(clk), .QN(
        \xmem_inst/mem[36][27] ) );
  DFF_X1 \xmem_inst/mem_reg[36][25]  ( .D(n5261), .CK(clk), .QN(
        \xmem_inst/mem[36][25] ) );
  DFF_X1 \xmem_inst/mem_reg[36][14]  ( .D(n5250), .CK(clk), .QN(
        \xmem_inst/mem[36][14] ) );
  DFF_X1 \xmem_inst/mem_reg[36][11]  ( .D(n5247), .CK(clk), .QN(
        \xmem_inst/mem[36][11] ) );
  DFF_X1 \xmem_inst/mem_reg[36][9]  ( .D(n5245), .CK(clk), .QN(
        \xmem_inst/mem[36][9] ) );
  DFF_X1 \xmem_inst/mem_reg[36][8]  ( .D(n5244), .CK(clk), .QN(
        \xmem_inst/mem[36][8] ) );
  DFF_X1 \xmem_inst/mem_reg[36][7]  ( .D(n5243), .CK(clk), .QN(
        \xmem_inst/mem[36][7] ) );
  DFF_X1 \xmem_inst/mem_reg[36][6]  ( .D(n5242), .CK(clk), .QN(
        \xmem_inst/mem[36][6] ) );
  DFF_X1 \xmem_inst/mem_reg[36][5]  ( .D(n5241), .CK(clk), .QN(
        \xmem_inst/mem[36][5] ) );
  DFF_X1 \xmem_inst/mem_reg[35][29]  ( .D(n5233), .CK(clk), .QN(
        \xmem_inst/mem[35][29] ) );
  DFF_X1 \xmem_inst/mem_reg[35][27]  ( .D(n5231), .CK(clk), .QN(
        \xmem_inst/mem[35][27] ) );
  DFF_X1 \xmem_inst/mem_reg[35][25]  ( .D(n5229), .CK(clk), .QN(
        \xmem_inst/mem[35][25] ) );
  DFF_X1 \xmem_inst/mem_reg[35][14]  ( .D(n5218), .CK(clk), .QN(
        \xmem_inst/mem[35][14] ) );
  DFF_X1 \xmem_inst/mem_reg[35][11]  ( .D(n5216), .CK(clk), .QN(
        \xmem_inst/mem[35][11] ) );
  DFF_X1 \xmem_inst/mem_reg[35][9]  ( .D(n5214), .CK(clk), .QN(
        \xmem_inst/mem[35][9] ) );
  DFF_X1 \xmem_inst/mem_reg[35][8]  ( .D(n5213), .CK(clk), .QN(
        \xmem_inst/mem[35][8] ) );
  DFF_X1 \xmem_inst/mem_reg[35][7]  ( .D(n5212), .CK(clk), .QN(
        \xmem_inst/mem[35][7] ) );
  DFF_X1 \xmem_inst/mem_reg[35][6]  ( .D(n5211), .CK(clk), .QN(
        \xmem_inst/mem[35][6] ) );
  DFF_X1 \xmem_inst/mem_reg[35][5]  ( .D(n5210), .CK(clk), .QN(
        \xmem_inst/mem[35][5] ) );
  DFF_X1 \xmem_inst/mem_reg[38][28]  ( .D(n5328), .CK(clk), .QN(
        \xmem_inst/mem[38][28] ) );
  DFF_X1 \xmem_inst/mem_reg[38][26]  ( .D(n5326), .CK(clk), .QN(
        \xmem_inst/mem[38][26] ) );
  DFF_X1 \xmem_inst/mem_reg[38][24]  ( .D(n5324), .CK(clk), .QN(
        \xmem_inst/mem[38][24] ) );
  DFF_X1 \xmem_inst/mem_reg[38][23]  ( .D(n5323), .CK(clk), .QN(
        \xmem_inst/mem[38][23] ) );
  DFF_X1 \xmem_inst/mem_reg[38][22]  ( .D(n5322), .CK(clk), .QN(
        \xmem_inst/mem[38][22] ) );
  DFF_X1 \xmem_inst/mem_reg[38][21]  ( .D(n5321), .CK(clk), .QN(
        \xmem_inst/mem[38][21] ) );
  DFF_X1 \xmem_inst/mem_reg[38][20]  ( .D(n5320), .CK(clk), .QN(
        \xmem_inst/mem[38][20] ) );
  DFF_X1 \xmem_inst/mem_reg[38][18]  ( .D(n5318), .CK(clk), .QN(
        \xmem_inst/mem[38][18] ) );
  DFF_X1 \xmem_inst/mem_reg[38][17]  ( .D(n5317), .CK(clk), .QN(
        \xmem_inst/mem[38][17] ) );
  DFF_X1 \xmem_inst/mem_reg[38][15]  ( .D(n5315), .CK(clk), .QN(
        \xmem_inst/mem[38][15] ) );
  DFF_X1 \xmem_inst/mem_reg[38][13]  ( .D(n5313), .CK(clk), .QN(
        \xmem_inst/mem[38][13] ) );
  DFF_X1 \xmem_inst/mem_reg[38][12]  ( .D(n5312), .CK(clk), .QN(
        \xmem_inst/mem[38][12] ) );
  DFF_X1 \xmem_inst/mem_reg[38][10]  ( .D(n5310), .CK(clk), .QN(
        \xmem_inst/mem[38][10] ) );
  DFF_X1 \xmem_inst/mem_reg[38][4]  ( .D(n5304), .CK(clk), .QN(
        \xmem_inst/mem[38][4] ) );
  DFF_X1 \xmem_inst/mem_reg[38][3]  ( .D(n5303), .CK(clk), .QN(
        \xmem_inst/mem[38][3] ) );
  DFF_X1 \xmem_inst/mem_reg[38][2]  ( .D(n5302), .CK(clk), .QN(
        \xmem_inst/mem[38][2] ) );
  DFF_X1 \xmem_inst/mem_reg[38][1]  ( .D(n5301), .CK(clk), .QN(
        \xmem_inst/mem[38][1] ) );
  DFF_X1 \xmem_inst/mem_reg[38][0]  ( .D(n5300), .CK(clk), .QN(
        \xmem_inst/mem[38][0] ) );
  DFF_X1 \xmem_inst/mem_reg[37][28]  ( .D(n5296), .CK(clk), .QN(
        \xmem_inst/mem[37][28] ) );
  DFF_X1 \xmem_inst/mem_reg[37][26]  ( .D(n5294), .CK(clk), .QN(
        \xmem_inst/mem[37][26] ) );
  DFF_X1 \xmem_inst/mem_reg[37][24]  ( .D(n5292), .CK(clk), .QN(
        \xmem_inst/mem[37][24] ) );
  DFF_X1 \xmem_inst/mem_reg[37][23]  ( .D(n5291), .CK(clk), .QN(
        \xmem_inst/mem[37][23] ) );
  DFF_X1 \xmem_inst/mem_reg[37][22]  ( .D(n5290), .CK(clk), .QN(
        \xmem_inst/mem[37][22] ) );
  DFF_X1 \xmem_inst/mem_reg[37][21]  ( .D(n5289), .CK(clk), .QN(
        \xmem_inst/mem[37][21] ) );
  DFF_X1 \xmem_inst/mem_reg[37][20]  ( .D(n5288), .CK(clk), .QN(
        \xmem_inst/mem[37][20] ) );
  DFF_X1 \xmem_inst/mem_reg[37][18]  ( .D(n5286), .CK(clk), .QN(
        \xmem_inst/mem[37][18] ) );
  DFF_X1 \xmem_inst/mem_reg[37][17]  ( .D(n5285), .CK(clk), .QN(
        \xmem_inst/mem[37][17] ) );
  DFF_X1 \xmem_inst/mem_reg[37][15]  ( .D(n5283), .CK(clk), .QN(
        \xmem_inst/mem[37][15] ) );
  DFF_X1 \xmem_inst/mem_reg[37][13]  ( .D(n5281), .CK(clk), .QN(
        \xmem_inst/mem[37][13] ) );
  DFF_X1 \xmem_inst/mem_reg[37][12]  ( .D(n5280), .CK(clk), .QN(
        \xmem_inst/mem[37][12] ) );
  DFF_X1 \xmem_inst/mem_reg[37][10]  ( .D(n5278), .CK(clk), .QN(
        \xmem_inst/mem[37][10] ) );
  DFF_X1 \xmem_inst/mem_reg[37][4]  ( .D(n5272), .CK(clk), .QN(
        \xmem_inst/mem[37][4] ) );
  DFF_X1 \xmem_inst/mem_reg[37][3]  ( .D(n5271), .CK(clk), .QN(
        \xmem_inst/mem[37][3] ) );
  DFF_X1 \xmem_inst/mem_reg[37][2]  ( .D(n5270), .CK(clk), .QN(
        \xmem_inst/mem[37][2] ) );
  DFF_X1 \xmem_inst/mem_reg[37][1]  ( .D(n5269), .CK(clk), .QN(
        \xmem_inst/mem[37][1] ) );
  DFF_X1 \xmem_inst/mem_reg[37][0]  ( .D(n5268), .CK(clk), .QN(
        \xmem_inst/mem[37][0] ) );
  DFF_X1 \xmem_inst/mem_reg[36][28]  ( .D(n5264), .CK(clk), .QN(
        \xmem_inst/mem[36][28] ) );
  DFF_X1 \xmem_inst/mem_reg[36][26]  ( .D(n5262), .CK(clk), .QN(
        \xmem_inst/mem[36][26] ) );
  DFF_X1 \xmem_inst/mem_reg[36][24]  ( .D(n5260), .CK(clk), .QN(
        \xmem_inst/mem[36][24] ) );
  DFF_X1 \xmem_inst/mem_reg[36][23]  ( .D(n5259), .CK(clk), .QN(
        \xmem_inst/mem[36][23] ) );
  DFF_X1 \xmem_inst/mem_reg[36][22]  ( .D(n5258), .CK(clk), .QN(
        \xmem_inst/mem[36][22] ) );
  DFF_X1 \xmem_inst/mem_reg[36][21]  ( .D(n5257), .CK(clk), .QN(
        \xmem_inst/mem[36][21] ) );
  DFF_X1 \xmem_inst/mem_reg[36][20]  ( .D(n5256), .CK(clk), .QN(
        \xmem_inst/mem[36][20] ) );
  DFF_X1 \xmem_inst/mem_reg[36][18]  ( .D(n5254), .CK(clk), .QN(
        \xmem_inst/mem[36][18] ) );
  DFF_X1 \xmem_inst/mem_reg[36][17]  ( .D(n5253), .CK(clk), .QN(
        \xmem_inst/mem[36][17] ) );
  DFF_X1 \xmem_inst/mem_reg[36][15]  ( .D(n5251), .CK(clk), .QN(
        \xmem_inst/mem[36][15] ) );
  DFF_X1 \xmem_inst/mem_reg[36][13]  ( .D(n5249), .CK(clk), .QN(
        \xmem_inst/mem[36][13] ) );
  DFF_X1 \xmem_inst/mem_reg[36][12]  ( .D(n5248), .CK(clk), .QN(
        \xmem_inst/mem[36][12] ) );
  DFF_X1 \xmem_inst/mem_reg[36][10]  ( .D(n5246), .CK(clk), .QN(
        \xmem_inst/mem[36][10] ) );
  DFF_X1 \xmem_inst/mem_reg[36][4]  ( .D(n5240), .CK(clk), .QN(
        \xmem_inst/mem[36][4] ) );
  DFF_X1 \xmem_inst/mem_reg[36][3]  ( .D(n5239), .CK(clk), .QN(
        \xmem_inst/mem[36][3] ) );
  DFF_X1 \xmem_inst/mem_reg[36][2]  ( .D(n5238), .CK(clk), .QN(
        \xmem_inst/mem[36][2] ) );
  DFF_X1 \xmem_inst/mem_reg[36][1]  ( .D(n5237), .CK(clk), .QN(
        \xmem_inst/mem[36][1] ) );
  DFF_X1 \xmem_inst/mem_reg[36][0]  ( .D(n5236), .CK(clk), .QN(
        \xmem_inst/mem[36][0] ) );
  DFF_X1 \xmem_inst/mem_reg[35][28]  ( .D(n5232), .CK(clk), .QN(
        \xmem_inst/mem[35][28] ) );
  DFF_X1 \xmem_inst/mem_reg[35][26]  ( .D(n5230), .CK(clk), .QN(
        \xmem_inst/mem[35][26] ) );
  DFF_X1 \xmem_inst/mem_reg[35][24]  ( .D(n5228), .CK(clk), .QN(
        \xmem_inst/mem[35][24] ) );
  DFF_X1 \xmem_inst/mem_reg[35][23]  ( .D(n5227), .CK(clk), .QN(
        \xmem_inst/mem[35][23] ) );
  DFF_X1 \xmem_inst/mem_reg[35][22]  ( .D(n5226), .CK(clk), .QN(
        \xmem_inst/mem[35][22] ) );
  DFF_X1 \xmem_inst/mem_reg[35][21]  ( .D(n5225), .CK(clk), .QN(
        \xmem_inst/mem[35][21] ) );
  DFF_X1 \xmem_inst/mem_reg[35][20]  ( .D(n5224), .CK(clk), .QN(
        \xmem_inst/mem[35][20] ) );
  DFF_X1 \xmem_inst/mem_reg[35][18]  ( .D(n5222), .CK(clk), .QN(
        \xmem_inst/mem[35][18] ) );
  DFF_X1 \xmem_inst/mem_reg[35][17]  ( .D(n5221), .CK(clk), .QN(
        \xmem_inst/mem[35][17] ) );
  DFF_X1 \xmem_inst/mem_reg[35][15]  ( .D(n5219), .CK(clk), .QN(
        \xmem_inst/mem[35][15] ) );
  DFF_X1 \xmem_inst/mem_reg[35][13]  ( .D(n5217), .CK(clk), .QN(
        \xmem_inst/mem[35][13] ) );
  DFF_X1 \xmem_inst/mem_reg[35][10]  ( .D(n5215), .CK(clk), .QN(
        \xmem_inst/mem[35][10] ) );
  DFF_X1 \xmem_inst/mem_reg[35][4]  ( .D(n5209), .CK(clk), .QN(
        \xmem_inst/mem[35][4] ) );
  DFF_X1 \xmem_inst/mem_reg[35][3]  ( .D(n5208), .CK(clk), .QN(
        \xmem_inst/mem[35][3] ) );
  DFF_X1 \xmem_inst/mem_reg[35][2]  ( .D(n5207), .CK(clk), .QN(
        \xmem_inst/mem[35][2] ) );
  DFF_X1 \xmem_inst/mem_reg[35][1]  ( .D(n5206), .CK(clk), .QN(
        \xmem_inst/mem[35][1] ) );
  DFF_X1 \xmem_inst/mem_reg[35][0]  ( .D(n5205), .CK(clk), .QN(
        \xmem_inst/mem[35][0] ) );
  DFF_X1 \xmem_inst/mem_reg[39][31]  ( .D(n5362), .CK(clk), .QN(
        \xmem_inst/mem[39][31] ) );
  DFF_X1 \xmem_inst/mem_reg[39][30]  ( .D(n5361), .CK(clk), .QN(
        \xmem_inst/mem[39][30] ) );
  DFF_X1 \xmem_inst/mem_reg[39][19]  ( .D(n5350), .CK(clk), .QN(
        \xmem_inst/mem[39][19] ) );
  DFF_X1 \xmem_inst/mem_reg[39][15]  ( .D(n5346), .CK(clk), .QN(
        \xmem_inst/mem[39][15] ) );
  DFF_X1 \xmem_inst/mem_reg[34][31]  ( .D(n5204), .CK(clk), .QN(
        \xmem_inst/mem[34][31] ) );
  DFF_X1 \xmem_inst/mem_reg[34][30]  ( .D(n5203), .CK(clk), .QN(
        \xmem_inst/mem[34][30] ) );
  DFF_X1 \xmem_inst/mem_reg[34][19]  ( .D(n5195), .CK(clk), .QN(
        \xmem_inst/mem[34][19] ) );
  DFF_X1 \xmem_inst/mem_reg[34][15]  ( .D(n5191), .CK(clk), .QN(
        \xmem_inst/mem[34][15] ) );
  DFF_X1 \xmem_inst/mem_reg[33][31]  ( .D(n5182), .CK(clk), .QN(
        \xmem_inst/mem[33][31] ) );
  DFF_X1 \xmem_inst/mem_reg[33][30]  ( .D(n5181), .CK(clk), .QN(
        \xmem_inst/mem[33][30] ) );
  DFF_X1 \xmem_inst/mem_reg[33][19]  ( .D(n5173), .CK(clk), .QN(
        \xmem_inst/mem[33][19] ) );
  DFF_X1 \xmem_inst/mem_reg[33][15]  ( .D(n5172), .CK(clk), .QN(
        \xmem_inst/mem[33][15] ) );
  DFF_X1 \xmem_inst/mem_reg[32][31]  ( .D(n5171), .CK(clk), .QN(
        \xmem_inst/mem[32][31] ) );
  DFF_X1 \xmem_inst/mem_reg[32][30]  ( .D(n5170), .CK(clk), .QN(
        \xmem_inst/mem[32][30] ) );
  DFF_X1 \xmem_inst/mem_reg[32][19]  ( .D(n5169), .CK(clk), .QN(
        \xmem_inst/mem[32][19] ) );
  DFF_X1 \xmem_inst/mem_reg[32][15]  ( .D(n5168), .CK(clk), .QN(
        \xmem_inst/mem[32][15] ) );
  DFF_X1 \xmem_inst/mem_reg[39][29]  ( .D(n5360), .CK(clk), .QN(
        \xmem_inst/mem[39][29] ) );
  DFF_X1 \xmem_inst/mem_reg[39][27]  ( .D(n5358), .CK(clk), .QN(
        \xmem_inst/mem[39][27] ) );
  DFF_X1 \xmem_inst/mem_reg[39][25]  ( .D(n5356), .CK(clk), .QN(
        \xmem_inst/mem[39][25] ) );
  DFF_X1 \xmem_inst/mem_reg[39][14]  ( .D(n5345), .CK(clk), .QN(
        \xmem_inst/mem[39][14] ) );
  DFF_X1 \xmem_inst/mem_reg[39][11]  ( .D(n5342), .CK(clk), .QN(
        \xmem_inst/mem[39][11] ) );
  DFF_X1 \xmem_inst/mem_reg[39][9]  ( .D(n5340), .CK(clk), .QN(
        \xmem_inst/mem[39][9] ) );
  DFF_X1 \xmem_inst/mem_reg[39][8]  ( .D(n5339), .CK(clk), .QN(
        \xmem_inst/mem[39][8] ) );
  DFF_X1 \xmem_inst/mem_reg[39][7]  ( .D(n5338), .CK(clk), .QN(
        \xmem_inst/mem[39][7] ) );
  DFF_X1 \xmem_inst/mem_reg[39][6]  ( .D(n5337), .CK(clk), .QN(
        \xmem_inst/mem[39][6] ) );
  DFF_X1 \xmem_inst/mem_reg[39][5]  ( .D(n5336), .CK(clk), .QN(
        \xmem_inst/mem[39][5] ) );
  DFF_X1 \xmem_inst/mem_reg[39][28]  ( .D(n5359), .CK(clk), .QN(
        \xmem_inst/mem[39][28] ) );
  DFF_X1 \xmem_inst/mem_reg[39][26]  ( .D(n5357), .CK(clk), .QN(
        \xmem_inst/mem[39][26] ) );
  DFF_X1 \xmem_inst/mem_reg[39][24]  ( .D(n5355), .CK(clk), .QN(
        \xmem_inst/mem[39][24] ) );
  DFF_X1 \xmem_inst/mem_reg[39][23]  ( .D(n5354), .CK(clk), .QN(
        \xmem_inst/mem[39][23] ) );
  DFF_X1 \xmem_inst/mem_reg[39][22]  ( .D(n5353), .CK(clk), .QN(
        \xmem_inst/mem[39][22] ) );
  DFF_X1 \xmem_inst/mem_reg[39][21]  ( .D(n5352), .CK(clk), .QN(
        \xmem_inst/mem[39][21] ) );
  DFF_X1 \xmem_inst/mem_reg[39][20]  ( .D(n5351), .CK(clk), .QN(
        \xmem_inst/mem[39][20] ) );
  DFF_X1 \xmem_inst/mem_reg[39][18]  ( .D(n5349), .CK(clk), .QN(
        \xmem_inst/mem[39][18] ) );
  DFF_X1 \xmem_inst/mem_reg[39][17]  ( .D(n5348), .CK(clk), .QN(
        \xmem_inst/mem[39][17] ) );
  DFF_X1 \xmem_inst/mem_reg[39][16]  ( .D(n5347), .CK(clk), .QN(
        \xmem_inst/mem[39][16] ) );
  DFF_X1 \xmem_inst/mem_reg[39][13]  ( .D(n5344), .CK(clk), .QN(
        \xmem_inst/mem[39][13] ) );
  DFF_X1 \xmem_inst/mem_reg[39][12]  ( .D(n5343), .CK(clk), .QN(
        \xmem_inst/mem[39][12] ) );
  DFF_X1 \xmem_inst/mem_reg[39][10]  ( .D(n5341), .CK(clk), .QN(
        \xmem_inst/mem[39][10] ) );
  DFF_X1 \xmem_inst/mem_reg[39][3]  ( .D(n5335), .CK(clk), .QN(
        \xmem_inst/mem[39][3] ) );
  DFF_X1 \xmem_inst/mem_reg[39][2]  ( .D(n5334), .CK(clk), .QN(
        \xmem_inst/mem[39][2] ) );
  DFF_X1 \xmem_inst/mem_reg[39][1]  ( .D(n5333), .CK(clk), .QN(
        \xmem_inst/mem[39][1] ) );
  DFF_X1 \xmem_inst/mem_reg[39][0]  ( .D(n5332), .CK(clk), .QN(
        \xmem_inst/mem[39][0] ) );
  DFF_X1 \xmem_inst/mem_reg[34][28]  ( .D(n5202), .CK(clk), .QN(
        \xmem_inst/mem[34][28] ) );
  DFF_X1 \xmem_inst/mem_reg[34][26]  ( .D(n5201), .CK(clk), .QN(
        \xmem_inst/mem[34][26] ) );
  DFF_X1 \xmem_inst/mem_reg[34][24]  ( .D(n5200), .CK(clk), .QN(
        \xmem_inst/mem[34][24] ) );
  DFF_X1 \xmem_inst/mem_reg[34][23]  ( .D(n5199), .CK(clk), .QN(
        \xmem_inst/mem[34][23] ) );
  DFF_X1 \xmem_inst/mem_reg[34][22]  ( .D(n5198), .CK(clk), .QN(
        \xmem_inst/mem[34][22] ) );
  DFF_X1 \xmem_inst/mem_reg[34][21]  ( .D(n5197), .CK(clk), .QN(
        \xmem_inst/mem[34][21] ) );
  DFF_X1 \xmem_inst/mem_reg[34][20]  ( .D(n5196), .CK(clk), .QN(
        \xmem_inst/mem[34][20] ) );
  DFF_X1 \xmem_inst/mem_reg[34][18]  ( .D(n5194), .CK(clk), .QN(
        \xmem_inst/mem[34][18] ) );
  DFF_X1 \xmem_inst/mem_reg[34][17]  ( .D(n5193), .CK(clk), .QN(
        \xmem_inst/mem[34][17] ) );
  DFF_X1 \xmem_inst/mem_reg[34][16]  ( .D(n5192), .CK(clk), .QN(
        \xmem_inst/mem[34][16] ) );
  DFF_X1 \xmem_inst/mem_reg[34][13]  ( .D(n5190), .CK(clk), .QN(
        \xmem_inst/mem[34][13] ) );
  DFF_X1 \xmem_inst/mem_reg[34][12]  ( .D(n5189), .CK(clk), .QN(
        \xmem_inst/mem[34][12] ) );
  DFF_X1 \xmem_inst/mem_reg[34][10]  ( .D(n5188), .CK(clk), .QN(
        \xmem_inst/mem[34][10] ) );
  DFF_X1 \xmem_inst/mem_reg[34][4]  ( .D(n5187), .CK(clk), .QN(
        \xmem_inst/mem[34][4] ) );
  DFF_X1 \xmem_inst/mem_reg[34][3]  ( .D(n5186), .CK(clk), .QN(
        \xmem_inst/mem[34][3] ) );
  DFF_X1 \xmem_inst/mem_reg[34][2]  ( .D(n5185), .CK(clk), .QN(
        \xmem_inst/mem[34][2] ) );
  DFF_X1 \xmem_inst/mem_reg[34][1]  ( .D(n5184), .CK(clk), .QN(
        \xmem_inst/mem[34][1] ) );
  DFF_X1 \xmem_inst/mem_reg[34][0]  ( .D(n5183), .CK(clk), .QN(
        \xmem_inst/mem[34][0] ) );
  DFF_X1 \xmem_inst/mem_reg[33][28]  ( .D(n5180), .CK(clk), .QN(
        \xmem_inst/mem[33][28] ) );
  DFF_X1 \xmem_inst/mem_reg[33][26]  ( .D(n5179), .CK(clk), .QN(
        \xmem_inst/mem[33][26] ) );
  DFF_X1 \xmem_inst/mem_reg[33][24]  ( .D(n5178), .CK(clk), .QN(
        \xmem_inst/mem[33][24] ) );
  DFF_X1 \xmem_inst/mem_reg[33][23]  ( .D(n5177), .CK(clk), .QN(
        \xmem_inst/mem[33][23] ) );
  DFF_X1 \xmem_inst/mem_reg[33][22]  ( .D(n5176), .CK(clk), .QN(
        \xmem_inst/mem[33][22] ) );
  DFF_X1 \xmem_inst/mem_reg[33][21]  ( .D(n5175), .CK(clk), .QN(
        \xmem_inst/mem[33][21] ) );
  DFF_X1 \xmem_inst/mem_reg[33][20]  ( .D(n5174), .CK(clk), .QN(
        \xmem_inst/mem[33][20] ) );
  SDFFS_X1 \fmem_inst/z_reg[0]  ( .D(\fmem_inst/N62 ), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(1'b1), .Q(fmem_data[0]), .QN(n283) );
  DFF_X2 \mac_unit_inst/adder_reg_reg[31]  ( .D(\mac_unit_inst/n81 ), .CK(clk), 
        .Q(\mac_unit_inst/adder_reg [31]), .QN(n309) );
  DFF_X2 \fmem_inst/z_reg[4]  ( .D(\fmem_inst/N66 ), .CK(clk), .Q(fmem_data[4]), .QN(n232) );
  DFF_X2 \fmem_inst/z_reg[15]  ( .D(\fmem_inst/N77 ), .CK(clk), .Q(
        fmem_data[15]), .QN(n282) );
  DFF_X2 \fmem_inst/z_reg[1]  ( .D(\fmem_inst/N63 ), .CK(clk), .Q(fmem_data[1]), .QN(n204) );
  DFF_X2 \fmem_inst/z_reg[14]  ( .D(\fmem_inst/N76 ), .CK(clk), .Q(
        fmem_data[14]), .QN(n280) );
  DFF_X2 \fmem_inst/z_reg[2]  ( .D(\fmem_inst/N64 ), .CK(clk), .Q(fmem_data[2]), .QN(n209) );
  DFF_X2 \fmem_inst/z_reg[6]  ( .D(\fmem_inst/N68 ), .CK(clk), .Q(fmem_data[6]), .QN(n4063) );
  DFF_X2 \xmem_inst/data_out_reg[0]  ( .D(\xmem_inst/N279 ), .CK(clk), .Q(
        xmem_data[0]), .QN(n315) );
  DFF_X1 \fmem_inst/z_reg[3]  ( .D(\fmem_inst/N65 ), .CK(clk), .Q(fmem_data[3]), .QN(n250) );
  DFF_X2 \mac_unit_inst/x_mult_f_reg_reg[19]  ( .D(\mac_unit_inst/n132 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [19]), .QN(n4143) );
  DFF_X2 \mac_unit_inst/x_mult_f_reg_reg[23]  ( .D(\mac_unit_inst/n136 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [23]), .QN(n4139) );
  DFF_X1 \fmem_inst/z_reg[10]  ( .D(\fmem_inst/N72 ), .CK(clk), .Q(
        fmem_data[10]), .QN(n202) );
  DFF_X1 \fmem_inst/z_reg[13]  ( .D(\fmem_inst/N75 ), .CK(clk), .Q(
        fmem_data[13]), .QN(n193) );
  DFF_X1 \fmem_inst/z_reg[7]  ( .D(\fmem_inst/N69 ), .CK(clk), .Q(fmem_data[7]), .QN(n262) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[24]  ( .D(\mac_unit_inst/n137 ), .CK(
        clk), .Q(\mac_unit_inst/x_mult_f_reg [24]), .QN(n4138) );
  XNOR2_X1 U148 ( .A(n1263), .B(n1261), .ZN(n132) );
  BUF_X1 U149 ( .A(n1731), .Z(n256) );
  NAND2_X1 U150 ( .A1(n131), .A2(n130), .ZN(n1285) );
  OAI21_X1 U151 ( .B1(n1262), .B2(n1263), .A(n1261), .ZN(n131) );
  BUF_X1 U152 ( .A(fmem_data[0]), .Z(n287) );
  NAND2_X2 U153 ( .A1(n406), .A2(n364), .ZN(n201) );
  BUF_X1 U154 ( .A(fmem_data[0]), .Z(n285) );
  INV_X1 U155 ( .A(n202), .ZN(n203) );
  BUF_X1 U156 ( .A(n2029), .Z(n185) );
  AOI21_X2 U157 ( .B1(n2033), .B2(n2032), .A(n2031), .ZN(n3552) );
  NAND2_X4 U158 ( .A1(n3291), .A2(n2604), .ZN(n2223) );
  NAND2_X1 U159 ( .A1(n122), .A2(n2203), .ZN(\mac_unit_inst/n122 ) );
  AOI21_X1 U160 ( .B1(n3657), .B2(n2170), .A(n2169), .ZN(n122) );
  NAND3_X1 U161 ( .A1(n123), .A2(n3658), .A3(n346), .ZN(\mac_unit_inst/n142 )
         );
  NAND2_X1 U162 ( .A1(n2072), .A2(n3680), .ZN(n123) );
  NAND2_X1 U163 ( .A1(n124), .A2(n2203), .ZN(\mac_unit_inst/n125 ) );
  AOI21_X1 U164 ( .B1(n3657), .B2(n2088), .A(n2087), .ZN(n124) );
  NAND2_X1 U165 ( .A1(n125), .A2(n2203), .ZN(\mac_unit_inst/n127 ) );
  AOI21_X1 U166 ( .B1(n3657), .B2(n2097), .A(n2096), .ZN(n125) );
  NAND2_X1 U167 ( .A1(n126), .A2(n2203), .ZN(\mac_unit_inst/n124 ) );
  AOI21_X1 U168 ( .B1(n3657), .B2(n2104), .A(n2103), .ZN(n126) );
  NAND2_X1 U169 ( .A1(n127), .A2(n2203), .ZN(\mac_unit_inst/n135 ) );
  AOI21_X1 U170 ( .B1(n3680), .B2(n2137), .A(n2136), .ZN(n127) );
  NAND2_X1 U171 ( .A1(n128), .A2(n2203), .ZN(\mac_unit_inst/n128 ) );
  AOI21_X1 U172 ( .B1(n3680), .B2(n2162), .A(n2161), .ZN(n128) );
  NAND2_X1 U173 ( .A1(n129), .A2(n2203), .ZN(\mac_unit_inst/n114 ) );
  AOI21_X1 U174 ( .B1(n3680), .B2(n2194), .A(n2193), .ZN(n129) );
  NAND2_X2 U175 ( .A1(n1262), .A2(n1263), .ZN(n130) );
  XNOR2_X1 U176 ( .A(n132), .B(n1262), .ZN(n1475) );
  NOR2_X1 U177 ( .A1(n1810), .A2(n1811), .ZN(n1814) );
  NAND2_X1 U178 ( .A1(n134), .A2(n133), .ZN(n1811) );
  INV_X1 U179 ( .A(n1900), .ZN(n133) );
  INV_X1 U180 ( .A(n288), .ZN(n134) );
  NAND2_X1 U181 ( .A1(n135), .A2(n3681), .ZN(\mac_unit_inst/n137 ) );
  AOI21_X1 U182 ( .B1(n3667), .B2(n3657), .A(n136), .ZN(n135) );
  NOR2_X1 U183 ( .A1(n2223), .A2(n4138), .ZN(n136) );
  BUF_X1 U184 ( .A(n1237), .Z(n199) );
  BUF_X1 U185 ( .A(n385), .Z(n1036) );
  AND2_X1 U186 ( .A1(n1081), .A2(n1080), .ZN(n217) );
  BUF_X1 U187 ( .A(n2025), .Z(n3681) );
  OAI21_X1 U188 ( .B1(n1070), .B2(n1069), .A(n164), .ZN(n163) );
  NAND2_X1 U189 ( .A1(n1070), .A2(n1069), .ZN(n162) );
  CLKBUF_X1 U190 ( .A(n2090), .Z(n186) );
  BUF_X1 U191 ( .A(n3488), .Z(n3486) );
  OR2_X1 U192 ( .A1(n1079), .A2(n1078), .ZN(n2075) );
  OR2_X1 U193 ( .A1(n1799), .A2(n1798), .ZN(n2047) );
  OR2_X1 U194 ( .A1(n1801), .A2(n1800), .ZN(n2051) );
  BUF_X1 U195 ( .A(n3488), .Z(n3422) );
  INV_X1 U196 ( .A(n181), .ZN(n2092) );
  NAND2_X1 U197 ( .A1(n1304), .A2(n1303), .ZN(n142) );
  NOR2_X1 U198 ( .A1(n1658), .A2(n1657), .ZN(n172) );
  NAND2_X1 U199 ( .A1(n1658), .A2(n1657), .ZN(n171) );
  BUF_X1 U200 ( .A(n3210), .Z(n3569) );
  BUF_X1 U201 ( .A(n3209), .Z(n3570) );
  BUF_X1 U202 ( .A(n3202), .Z(n3604) );
  BUF_X1 U203 ( .A(n3147), .Z(n3572) );
  BUF_X1 U204 ( .A(n3148), .Z(n3602) );
  BUF_X1 U205 ( .A(n3598), .Z(n3233) );
  BUF_X1 U206 ( .A(n3251), .Z(n3584) );
  BUF_X1 U207 ( .A(n3189), .Z(n3571) );
  BUF_X1 U208 ( .A(n3573), .Z(n3244) );
  BUF_X1 U209 ( .A(n3084), .Z(n3585) );
  BUF_X1 U210 ( .A(n3586), .Z(n3253) );
  BUF_X1 U211 ( .A(n3591), .Z(n3179) );
  NAND2_X1 U212 ( .A1(n648), .A2(n647), .ZN(n175) );
  BUF_X1 U213 ( .A(n3599), .Z(n3226) );
  BUF_X1 U214 ( .A(n3184), .Z(n3613) );
  BUF_X1 U215 ( .A(n3203), .Z(n3580) );
  BUF_X1 U216 ( .A(n3153), .Z(n3568) );
  BUF_X1 U217 ( .A(n3250), .Z(n3574) );
  BUF_X1 U218 ( .A(n3178), .Z(n3630) );
  BUF_X1 U219 ( .A(n3072), .Z(n3629) );
  BUF_X1 U220 ( .A(n2967), .Z(n3614) );
  BUF_X1 U221 ( .A(n3618), .Z(n3252) );
  BUF_X1 U222 ( .A(n3154), .Z(n3616) );
  BUF_X1 U223 ( .A(n3254), .Z(n3624) );
  BUF_X1 U224 ( .A(n3234), .Z(n3615) );
  CLKBUF_X2 U225 ( .A(n1371), .Z(n296) );
  CLKBUF_X2 U226 ( .A(n383), .Z(n858) );
  CLKBUF_X2 U227 ( .A(n383), .Z(n801) );
  CLKBUF_X1 U228 ( .A(n1575), .Z(n244) );
  CLKBUF_X2 U229 ( .A(n357), .Z(n547) );
  CLKBUF_X2 U230 ( .A(n375), .Z(n1249) );
  BUF_X2 U231 ( .A(n373), .Z(n138) );
  BUF_X1 U232 ( .A(n249), .Z(n247) );
  BUF_X1 U233 ( .A(n1575), .Z(n245) );
  BUF_X1 U234 ( .A(fmem_data[3]), .Z(n228) );
  BUF_X1 U235 ( .A(xmem_data[15]), .Z(n1113) );
  BUF_X1 U236 ( .A(fmem_data[3]), .Z(n229) );
  CLKBUF_X2 U237 ( .A(xmem_data[5]), .Z(n791) );
  BUF_X1 U238 ( .A(xmem_data[1]), .Z(n225) );
  BUF_X2 U239 ( .A(xmem_data[5]), .Z(n261) );
  CLKBUF_X1 U240 ( .A(n329), .Z(n198) );
  BUF_X1 U241 ( .A(xmem_data[1]), .Z(n226) );
  CLKBUF_X1 U242 ( .A(n4062), .Z(n213) );
  BUF_X1 U243 ( .A(n2131), .Z(n218) );
  NAND2_X1 U244 ( .A1(n748), .A2(n747), .ZN(n2124) );
  OR2_X1 U245 ( .A1(n1984), .A2(n1983), .ZN(n1986) );
  CLKBUF_X1 U246 ( .A(n2028), .Z(n1859) );
  OR2_X1 U247 ( .A1(n1876), .A2(n1875), .ZN(n2042) );
  OR2_X1 U248 ( .A1(n1865), .A2(n1864), .ZN(n2149) );
  NOR2_X1 U249 ( .A1(n753), .A2(n752), .ZN(n1846) );
  INV_X1 U250 ( .A(n2076), .ZN(n139) );
  AOI21_X1 U251 ( .B1(n1838), .B2(n3650), .A(n1837), .ZN(n2183) );
  NOR2_X1 U252 ( .A1(n3296), .A2(n3295), .ZN(n3488) );
  NAND2_X1 U253 ( .A1(n1487), .A2(n1486), .ZN(n1877) );
  NAND2_X1 U254 ( .A1(n163), .A2(n162), .ZN(n1078) );
  OR2_X1 U255 ( .A1(n1994), .A2(n1995), .ZN(n1997) );
  NAND2_X1 U256 ( .A1(n1291), .A2(n1290), .ZN(n3555) );
  XNOR2_X1 U257 ( .A(n155), .B(n1480), .ZN(n1878) );
  NAND2_X1 U258 ( .A1(n1482), .A2(n1481), .ZN(n150) );
  NAND2_X1 U259 ( .A1(n143), .A2(n142), .ZN(n1345) );
  XNOR2_X1 U260 ( .A(n1482), .B(n1481), .ZN(n155) );
  OAI21_X1 U261 ( .B1(n1556), .B2(n1555), .A(n1554), .ZN(n1907) );
  OAI21_X1 U262 ( .B1(n1304), .B2(n1303), .A(n1302), .ZN(n143) );
  NOR2_X1 U263 ( .A1(n2002), .A2(n2001), .ZN(n1689) );
  NOR2_X1 U264 ( .A1(n589), .A2(n588), .ZN(n2179) );
  CLKBUF_X1 U265 ( .A(n433), .Z(n386) );
  OAI21_X1 U266 ( .B1(n173), .B2(n172), .A(n171), .ZN(n1688) );
  XNOR2_X1 U267 ( .A(n174), .B(n1656), .ZN(n1669) );
  XNOR2_X1 U268 ( .A(n1658), .B(n1657), .ZN(n174) );
  INV_X1 U269 ( .A(n1656), .ZN(n173) );
  XNOR2_X1 U270 ( .A(n149), .B(n462), .ZN(n598) );
  NAND2_X1 U271 ( .A1(n176), .A2(n175), .ZN(n733) );
  CLKBUF_X1 U272 ( .A(n3754), .Z(n3755) );
  CLKBUF_X1 U273 ( .A(n3719), .Z(n3720) );
  CLKBUF_X1 U274 ( .A(n3715), .Z(n3716) );
  OAI21_X1 U275 ( .B1(n648), .B2(n647), .A(n178), .ZN(n176) );
  CLKBUF_X1 U276 ( .A(n3711), .Z(n3712) );
  CLKBUF_X1 U277 ( .A(n4000), .Z(n4003) );
  CLKBUF_X1 U278 ( .A(n3707), .Z(n3708) );
  CLKBUF_X1 U279 ( .A(n3704), .Z(n3705) );
  CLKBUF_X1 U280 ( .A(n3701), .Z(n3702) );
  CLKBUF_X1 U281 ( .A(n3698), .Z(n3699) );
  CLKBUF_X1 U282 ( .A(n3776), .Z(n3777) );
  CLKBUF_X1 U283 ( .A(n3769), .Z(n3770) );
  CLKBUF_X1 U284 ( .A(n3766), .Z(n3767) );
  CLKBUF_X1 U285 ( .A(n3763), .Z(n3764) );
  CLKBUF_X1 U286 ( .A(n3760), .Z(n3761) );
  CLKBUF_X1 U287 ( .A(n3757), .Z(n3758) );
  CLKBUF_X1 U288 ( .A(n3856), .Z(n3858) );
  CLKBUF_X1 U289 ( .A(n3786), .Z(n3787) );
  CLKBUF_X1 U290 ( .A(n3741), .Z(n3742) );
  CLKBUF_X1 U291 ( .A(n3744), .Z(n3745) );
  NAND2_X1 U292 ( .A1(n462), .A2(n463), .ZN(n147) );
  CLKBUF_X1 U293 ( .A(n3747), .Z(n3748) );
  CLKBUF_X1 U294 ( .A(n2223), .Z(n3659) );
  CLKBUF_X1 U295 ( .A(n3802), .Z(n3803) );
  CLKBUF_X1 U296 ( .A(n3792), .Z(n3793) );
  CLKBUF_X1 U297 ( .A(n3795), .Z(n3796) );
  CLKBUF_X1 U298 ( .A(n3879), .Z(n3880) );
  CLKBUF_X1 U299 ( .A(n3751), .Z(n3752) );
  CLKBUF_X1 U300 ( .A(n3883), .Z(n3884) );
  CLKBUF_X1 U301 ( .A(n3798), .Z(n3799) );
  CLKBUF_X1 U302 ( .A(n3738), .Z(n3739) );
  CLKBUF_X1 U303 ( .A(n3887), .Z(n3888) );
  CLKBUF_X1 U304 ( .A(n3832), .Z(n3834) );
  CLKBUF_X1 U305 ( .A(n3725), .Z(n3726) );
  CLKBUF_X1 U306 ( .A(n3783), .Z(n3784) );
  CLKBUF_X1 U307 ( .A(n3963), .Z(n3966) );
  CLKBUF_X1 U308 ( .A(n3729), .Z(n3730) );
  CLKBUF_X1 U309 ( .A(n3732), .Z(n3733) );
  XNOR2_X1 U310 ( .A(n463), .B(n461), .ZN(n149) );
  CLKBUF_X1 U311 ( .A(n3927), .Z(n3930) );
  CLKBUF_X1 U312 ( .A(n3893), .Z(n3894) );
  CLKBUF_X1 U313 ( .A(n3876), .Z(n3877) );
  CLKBUF_X1 U314 ( .A(n3735), .Z(n3736) );
  CLKBUF_X1 U315 ( .A(n3869), .Z(n3871) );
  CLKBUF_X1 U316 ( .A(n3780), .Z(n3781) );
  CLKBUF_X1 U317 ( .A(n3789), .Z(n3790) );
  CLKBUF_X1 U318 ( .A(n3772), .Z(n3773) );
  BUF_X1 U319 ( .A(n2958), .Z(n3631) );
  BUF_X1 U320 ( .A(n3235), .Z(n3625) );
  CLKBUF_X1 U321 ( .A(n1371), .Z(n295) );
  BUF_X1 U322 ( .A(n1371), .Z(n297) );
  NAND4_X1 U323 ( .A1(xmem_addr[5]), .A2(n3896), .A3(n4083), .A4(n4081), .ZN(
        n3890) );
  NAND3_X1 U324 ( .A1(n3728), .A2(n3896), .A3(n4083), .ZN(n3723) );
  BUF_X1 U325 ( .A(n788), .Z(n1353) );
  CLKBUF_X2 U326 ( .A(n1575), .Z(n182) );
  CLKBUF_X2 U327 ( .A(n375), .Z(n1233) );
  XNOR2_X1 U328 ( .A(n228), .B(n281), .ZN(n1156) );
  BUF_X2 U329 ( .A(n352), .Z(n774) );
  BUF_X1 U330 ( .A(n230), .Z(n1271) );
  BUF_X1 U331 ( .A(n248), .Z(n1253) );
  BUF_X2 U332 ( .A(n207), .Z(n1641) );
  BUF_X1 U333 ( .A(n215), .Z(n191) );
  BUF_X1 U334 ( .A(n1096), .Z(n1638) );
  CLKBUF_X2 U335 ( .A(xmem_data[11]), .Z(n886) );
  INV_X1 U336 ( .A(n193), .ZN(n194) );
  BUF_X2 U337 ( .A(n215), .Z(n140) );
  BUF_X2 U338 ( .A(n230), .Z(n141) );
  BUF_X2 U339 ( .A(fmem_data[0]), .Z(n286) );
  INV_X1 U340 ( .A(n283), .ZN(n284) );
  INV_X1 U341 ( .A(n262), .ZN(n238) );
  CLKBUF_X1 U342 ( .A(fmem_data[3]), .Z(n227) );
  INV_X1 U343 ( .A(n280), .ZN(n188) );
  CLKBUF_X1 U344 ( .A(n4061), .Z(n214) );
  INV_X1 U345 ( .A(n282), .ZN(n192) );
  CLKBUF_X1 U346 ( .A(xmem_data[1]), .Z(n639) );
  INV_X1 U347 ( .A(n4057), .ZN(n184) );
  INV_X1 U348 ( .A(n257), .ZN(n258) );
  XNOR2_X1 U349 ( .A(n144), .B(n1302), .ZN(n1346) );
  XNOR2_X1 U350 ( .A(n1304), .B(n1303), .ZN(n144) );
  NAND2_X1 U351 ( .A1(n145), .A2(n3681), .ZN(\mac_unit_inst/n132 ) );
  AOI21_X1 U352 ( .B1(n3680), .B2(n3679), .A(n146), .ZN(n145) );
  NOR2_X1 U353 ( .A1(n2223), .A2(n4143), .ZN(n146) );
  NAND2_X1 U354 ( .A1(n2156), .A2(n2158), .ZN(n1845) );
  NOR2_X1 U355 ( .A1(n1842), .A2(n1828), .ZN(n2156) );
  NAND2_X1 U356 ( .A1(n148), .A2(n147), .ZN(n453) );
  OAI21_X1 U357 ( .B1(n462), .B2(n463), .A(n461), .ZN(n148) );
  NAND2_X1 U358 ( .A1(n151), .A2(n150), .ZN(n1875) );
  NAND2_X1 U359 ( .A1(n1480), .A2(n152), .ZN(n151) );
  NAND2_X1 U360 ( .A1(n154), .A2(n153), .ZN(n152) );
  INV_X1 U361 ( .A(n1481), .ZN(n153) );
  INV_X1 U362 ( .A(n1482), .ZN(n154) );
  NAND2_X1 U363 ( .A1(n3658), .A2(n156), .ZN(\mac_unit_inst/n126 ) );
  AOI21_X1 U364 ( .B1(n3657), .B2(n3649), .A(n157), .ZN(n156) );
  NOR2_X1 U365 ( .A1(n3659), .A2(n4125), .ZN(n157) );
  NAND2_X1 U366 ( .A1(n3658), .A2(n158), .ZN(\mac_unit_inst/n121 ) );
  AOI21_X1 U367 ( .B1(n3680), .B2(n3656), .A(n159), .ZN(n158) );
  NOR2_X1 U368 ( .A1(n3659), .A2(n4130), .ZN(n159) );
  NAND2_X1 U369 ( .A1(n160), .A2(n3681), .ZN(\mac_unit_inst/n129 ) );
  AOI21_X1 U370 ( .B1(n3657), .B2(n3644), .A(n161), .ZN(n160) );
  NOR2_X1 U371 ( .A1(n3659), .A2(n4122), .ZN(n161) );
  XNOR2_X1 U372 ( .A(xmem_data[15]), .B(n333), .ZN(n364) );
  XNOR2_X1 U373 ( .A(xmem_data[13]), .B(xmem_data[14]), .ZN(n406) );
  XNOR2_X1 U374 ( .A(n165), .B(n164), .ZN(n1865) );
  XNOR2_X1 U375 ( .A(n820), .B(n1059), .ZN(n164) );
  XNOR2_X1 U376 ( .A(n1070), .B(n1069), .ZN(n165) );
  BUF_X4 U377 ( .A(xmem_data[15]), .Z(n1269) );
  BUF_X4 U378 ( .A(n1123), .Z(n1743) );
  AND2_X1 U379 ( .A1(n1135), .A2(n166), .ZN(n168) );
  INV_X1 U380 ( .A(n1299), .ZN(n166) );
  OAI21_X1 U381 ( .B1(n168), .B2(n167), .A(n1136), .ZN(n1213) );
  INV_X1 U382 ( .A(n1301), .ZN(n167) );
  NAND2_X1 U383 ( .A1(n1138), .A2(n1137), .ZN(n1339) );
  NAND2_X1 U384 ( .A1(n1210), .A2(n1211), .ZN(n1137) );
  OAI21_X1 U385 ( .B1(n1210), .B2(n1211), .A(n1213), .ZN(n1138) );
  AOI21_X1 U386 ( .B1(n170), .B2(n169), .A(n2006), .ZN(n1936) );
  INV_X1 U387 ( .A(n1999), .ZN(n169) );
  INV_X1 U388 ( .A(n2000), .ZN(n170) );
  OAI21_X1 U389 ( .B1(n1853), .B2(n139), .A(n2132), .ZN(n1854) );
  AND2_X1 U390 ( .A1(n1079), .A2(n1078), .ZN(n2076) );
  XNOR2_X1 U391 ( .A(n177), .B(n648), .ZN(n689) );
  XNOR2_X1 U392 ( .A(n647), .B(n178), .ZN(n177) );
  OAI21_X1 U393 ( .B1(n641), .B2(n315), .A(n179), .ZN(n178) );
  OR2_X1 U394 ( .A1(n642), .A2(n640), .ZN(n179) );
  BUF_X1 U395 ( .A(n4059), .Z(n180) );
  AND2_X1 U396 ( .A1(n622), .A2(n621), .ZN(n181) );
  INV_X1 U397 ( .A(n273), .ZN(n183) );
  BUF_X1 U398 ( .A(n1127), .Z(n1732) );
  AND2_X1 U399 ( .A1(n1291), .A2(n1290), .ZN(n187) );
  INV_X1 U400 ( .A(n4051), .ZN(n189) );
  INV_X1 U401 ( .A(n189), .ZN(n190) );
  INV_X1 U402 ( .A(n217), .ZN(n2132) );
  XOR2_X1 U403 ( .A(n209), .B(n246), .Z(n1257) );
  BUF_X1 U404 ( .A(n899), .Z(n1532) );
  INV_X1 U405 ( .A(n1027), .ZN(n195) );
  BUF_X1 U406 ( .A(n1680), .Z(n196) );
  BUF_X1 U407 ( .A(n842), .Z(n197) );
  BUF_X2 U408 ( .A(n1255), .Z(n1237) );
  NAND2_X1 U409 ( .A1(n1148), .A2(n1147), .ZN(n200) );
  XOR2_X1 U410 ( .A(n204), .B(n244), .Z(n1238) );
  INV_X1 U411 ( .A(n1235), .ZN(n306) );
  INV_X1 U412 ( .A(n330), .ZN(n205) );
  INV_X1 U413 ( .A(n205), .ZN(n206) );
  XNOR2_X1 U414 ( .A(n330), .B(n221), .ZN(n207) );
  BUF_X1 U415 ( .A(n1869), .Z(n208) );
  XOR2_X1 U416 ( .A(n209), .B(n1324), .Z(n878) );
  INV_X1 U417 ( .A(n1874), .ZN(n210) );
  AND2_X1 U418 ( .A1(n1865), .A2(n1864), .ZN(n211) );
  XNOR2_X1 U419 ( .A(n212), .B(n339), .ZN(n352) );
  BUF_X1 U420 ( .A(n393), .Z(n931) );
  BUF_X4 U421 ( .A(n393), .Z(n1037) );
  XNOR2_X1 U422 ( .A(n4062), .B(n313), .ZN(n215) );
  NOR2_X2 U423 ( .A1(n587), .A2(n586), .ZN(n2164) );
  BUF_X4 U424 ( .A(n378), .Z(n871) );
  FA_X1 U425 ( .A(n1671), .B(n1670), .CI(n1669), .CO(n137), .S(n216) );
  AOI21_X1 U426 ( .B1(n1872), .B2(n1852), .A(n1855), .ZN(n2131) );
  BUF_X1 U427 ( .A(n230), .Z(n219) );
  XNOR2_X1 U428 ( .A(xmem_data[26]), .B(n312), .ZN(n1095) );
  BUF_X1 U429 ( .A(xmem_data[27]), .Z(n1096) );
  XNOR2_X1 U430 ( .A(n1900), .B(n220), .ZN(n1965) );
  XOR2_X1 U431 ( .A(n1184), .B(n259), .Z(n220) );
  XNOR2_X1 U432 ( .A(n330), .B(n221), .ZN(n852) );
  NOR2_X1 U433 ( .A1(n1885), .A2(n2026), .ZN(n222) );
  XNOR2_X1 U434 ( .A(xmem_data[17]), .B(n269), .ZN(n681) );
  XNOR2_X1 U435 ( .A(n4058), .B(n223), .ZN(n362) );
  XNOR2_X1 U436 ( .A(n4050), .B(n4051), .ZN(n224) );
  XNOR2_X1 U437 ( .A(xmem_data[14]), .B(xmem_data[13]), .ZN(n230) );
  BUF_X2 U438 ( .A(n1680), .Z(n274) );
  BUF_X1 U439 ( .A(n1123), .Z(n231) );
  INV_X1 U440 ( .A(n232), .ZN(n233) );
  BUF_X1 U441 ( .A(n1571), .Z(n234) );
  BUF_X1 U442 ( .A(n1571), .Z(n235) );
  CLKBUF_X1 U443 ( .A(n900), .Z(n1533) );
  XNOR2_X1 U444 ( .A(xmem_data[18]), .B(n4064), .ZN(n763) );
  OR2_X1 U445 ( .A1(n842), .A2(n841), .ZN(n236) );
  NOR2_X1 U446 ( .A1(n624), .A2(n623), .ZN(n237) );
  NOR2_X1 U447 ( .A1(n624), .A2(n623), .ZN(n1829) );
  OAI22_X1 U448 ( .A1(n1713), .A2(n1156), .B1(n1155), .B2(n1731), .ZN(n239) );
  BUF_X2 U449 ( .A(n402), .Z(n1251) );
  XOR2_X1 U450 ( .A(n825), .B(n826), .Z(n240) );
  XOR2_X1 U451 ( .A(n824), .B(n240), .Z(n831) );
  NAND2_X1 U452 ( .A1(n824), .A2(n825), .ZN(n241) );
  NAND2_X1 U453 ( .A1(n824), .A2(n826), .ZN(n242) );
  NAND2_X1 U454 ( .A1(n825), .A2(n826), .ZN(n243) );
  NAND3_X1 U455 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n1059) );
  XNOR2_X1 U456 ( .A(xmem_data[2]), .B(n329), .ZN(n351) );
  BUF_X2 U457 ( .A(xmem_data[25]), .Z(n246) );
  INV_X1 U458 ( .A(n4065), .ZN(n1575) );
  XNOR2_X1 U459 ( .A(n4059), .B(n4060), .ZN(n248) );
  XNOR2_X1 U460 ( .A(n4059), .B(n4060), .ZN(n249) );
  XNOR2_X1 U461 ( .A(n250), .B(n300), .ZN(n876) );
  NOR2_X1 U462 ( .A1(n1342), .A2(n299), .ZN(n251) );
  BUF_X4 U463 ( .A(xmem_data[13]), .Z(n252) );
  BUF_X2 U464 ( .A(xmem_data[13]), .Z(n1245) );
  NAND2_X1 U465 ( .A1(n1138), .A2(n1137), .ZN(n253) );
  BUF_X1 U466 ( .A(n1680), .Z(n275) );
  NOR3_X1 U467 ( .A1(n1750), .A2(n1791), .A3(n1749), .ZN(n254) );
  NOR3_X1 U468 ( .A1(n1750), .A2(n1791), .A3(n1749), .ZN(n1821) );
  BUF_X1 U469 ( .A(n1947), .Z(n255) );
  BUF_X1 U470 ( .A(n1337), .Z(n259) );
  OR2_X1 U471 ( .A1(n1008), .A2(n1120), .ZN(n260) );
  NAND2_X1 U472 ( .A1(n260), .A2(n1119), .ZN(n1172) );
  XNOR2_X1 U473 ( .A(n262), .B(n312), .ZN(n1311) );
  BUF_X4 U474 ( .A(n423), .Z(n1010) );
  BUF_X1 U475 ( .A(n373), .Z(n711) );
  AND2_X1 U476 ( .A1(n842), .A2(n841), .ZN(n263) );
  AND2_X1 U477 ( .A1(n1953), .A2(n1978), .ZN(n264) );
  XNOR2_X1 U478 ( .A(n4056), .B(n329), .ZN(n409) );
  BUF_X1 U479 ( .A(n1948), .Z(n265) );
  XNOR2_X1 U480 ( .A(n266), .B(n4068), .ZN(n363) );
  XNOR2_X1 U481 ( .A(n651), .B(n267), .ZN(n690) );
  XNOR2_X1 U482 ( .A(n650), .B(n649), .ZN(n267) );
  XNOR2_X1 U483 ( .A(n1950), .B(n1949), .ZN(n1951) );
  XNOR2_X1 U484 ( .A(n4058), .B(xmem_data[10]), .ZN(n347) );
  INV_X1 U485 ( .A(n1882), .ZN(n268) );
  OR2_X2 U486 ( .A1(n1081), .A2(n1080), .ZN(n2133) );
  XNOR2_X1 U487 ( .A(n269), .B(n4053), .ZN(n788) );
  XNOR2_X1 U488 ( .A(n270), .B(n4068), .ZN(n385) );
  XNOR2_X1 U489 ( .A(n271), .B(n198), .ZN(n401) );
  XNOR2_X1 U490 ( .A(xmem_data[29]), .B(n272), .ZN(n1101) );
  XNOR2_X1 U491 ( .A(n273), .B(n312), .ZN(n1159) );
  BUF_X2 U492 ( .A(n1680), .Z(n276) );
  NAND2_X1 U493 ( .A1(n1025), .A2(n1032), .ZN(n1680) );
  BUF_X2 U494 ( .A(n1127), .Z(n1713) );
  BUF_X4 U495 ( .A(n360), .Z(n857) );
  BUF_X1 U496 ( .A(n735), .Z(n277) );
  NAND3_X1 U497 ( .A1(n1954), .A2(n1955), .A3(n264), .ZN(n2017) );
  FA_X1 U498 ( .A(n1688), .B(n1687), .CI(n1686), .S(n278) );
  BUF_X4 U499 ( .A(xmem_data[7]), .Z(n279) );
  BUF_X2 U500 ( .A(xmem_data[7]), .Z(n849) );
  XOR2_X1 U501 ( .A(fmem_data[7]), .B(n206), .Z(n1275) );
  NAND2_X2 U502 ( .A1(n844), .A2(n852), .ZN(n1008) );
  XNOR2_X1 U503 ( .A(n4062), .B(n313), .ZN(n1032) );
  XNOR2_X1 U504 ( .A(xmem_data[12]), .B(n4061), .ZN(n361) );
  BUF_X2 U505 ( .A(xmem_data[29]), .Z(n1711) );
  XNOR2_X1 U506 ( .A(n280), .B(n4061), .ZN(n1250) );
  XOR2_X1 U507 ( .A(fmem_data[8]), .B(n206), .Z(n1197) );
  INV_X2 U508 ( .A(n331), .ZN(n281) );
  XNOR2_X1 U509 ( .A(n282), .B(n4061), .ZN(n1248) );
  XNOR2_X1 U510 ( .A(n1184), .B(n259), .ZN(n288) );
  NAND2_X1 U511 ( .A1(n651), .A2(n650), .ZN(n289) );
  NAND2_X1 U512 ( .A1(n651), .A2(n649), .ZN(n290) );
  NAND2_X1 U513 ( .A1(n650), .A2(n649), .ZN(n291) );
  NAND3_X1 U514 ( .A1(n289), .A2(n290), .A3(n291), .ZN(n734) );
  OAI211_X1 U515 ( .C1(n1826), .C2(n1825), .A(n1823), .B(n1824), .ZN(n292) );
  OAI211_X1 U516 ( .C1(n1826), .C2(n1825), .A(n1823), .B(n1824), .ZN(n3561) );
  AND2_X1 U517 ( .A1(n1797), .A2(n1796), .ZN(n293) );
  INV_X1 U518 ( .A(n1848), .ZN(n294) );
  NAND2_X1 U519 ( .A1(n347), .A2(n224), .ZN(n1371) );
  AOI21_X1 U520 ( .B1(n2076), .B2(n2133), .A(n217), .ZN(n298) );
  NOR2_X1 U521 ( .A1(n1811), .A2(n1810), .ZN(n299) );
  BUF_X2 U522 ( .A(n4064), .Z(n300) );
  OR2_X1 U523 ( .A1(n1878), .A2(n1877), .ZN(n301) );
  NAND2_X1 U524 ( .A1(n301), .A2(n2042), .ZN(n1885) );
  OAI21_X1 U525 ( .B1(n2147), .B2(n1858), .A(n1857), .ZN(n302) );
  AOI21_X1 U526 ( .B1(n2120), .B2(n1851), .A(n1850), .ZN(n303) );
  OAI21_X1 U527 ( .B1(n303), .B2(n1858), .A(n1857), .ZN(n3661) );
  BUF_X1 U528 ( .A(n3565), .Z(n304) );
  INV_X1 U529 ( .A(n306), .ZN(n305) );
  INV_X1 U530 ( .A(n1235), .ZN(n307) );
  INV_X1 U531 ( .A(n1235), .ZN(n1696) );
  NAND2_X1 U532 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U533 ( .A1(n1582), .A2(n1581), .ZN(n1608) );
  NAND2_X1 U534 ( .A1(n1178), .A2(n1177), .ZN(n1147) );
  OR2_X1 U535 ( .A1(n1178), .A2(n1177), .ZN(n1146) );
  NAND2_X1 U536 ( .A1(n1540), .A2(n1539), .ZN(n1569) );
  NAND2_X1 U537 ( .A1(n1566), .A2(n1565), .ZN(n1909) );
  OAI21_X1 U538 ( .B1(n1907), .B2(n1564), .A(n1563), .ZN(n1566) );
  NAND2_X1 U539 ( .A1(n1907), .A2(n1564), .ZN(n1565) );
  XNOR2_X1 U540 ( .A(n1523), .B(n1514), .ZN(n1553) );
  XNOR2_X1 U541 ( .A(n1525), .B(n1524), .ZN(n1514) );
  XNOR2_X1 U542 ( .A(n1415), .B(n1414), .ZN(n1400) );
  BUF_X2 U543 ( .A(n385), .Z(n929) );
  NAND2_X1 U544 ( .A1(n1341), .A2(n1340), .ZN(n1945) );
  NAND2_X1 U545 ( .A1(n253), .A2(n1338), .ZN(n1340) );
  OAI21_X1 U546 ( .B1(n1338), .B2(n253), .A(n1337), .ZN(n1341) );
  OAI21_X1 U547 ( .B1(n1384), .B2(n1383), .A(n1382), .ZN(n1437) );
  NAND2_X1 U548 ( .A1(n1431), .A2(n1430), .ZN(n1382) );
  OAI21_X1 U549 ( .B1(n1019), .B2(n1018), .A(n1017), .ZN(n1385) );
  NOR2_X1 U550 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  NAND2_X1 U551 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  INV_X1 U552 ( .A(n1049), .ZN(n1045) );
  XNOR2_X1 U553 ( .A(n1062), .B(n1061), .ZN(n1063) );
  INV_X1 U554 ( .A(n743), .ZN(n740) );
  XNOR2_X1 U555 ( .A(n705), .B(n684), .ZN(n743) );
  XNOR2_X1 U556 ( .A(n703), .B(n702), .ZN(n684) );
  INV_X1 U557 ( .A(n1874), .ZN(n2027) );
  XNOR2_X1 U558 ( .A(n938), .B(n999), .ZN(n1048) );
  OAI21_X1 U559 ( .B1(n1065), .B2(n1066), .A(n1067), .ZN(n987) );
  NAND2_X1 U560 ( .A1(n1066), .A2(n1065), .ZN(n986) );
  NAND2_X1 U561 ( .A1(n1062), .A2(n1061), .ZN(n963) );
  OR2_X1 U562 ( .A1(n1062), .A2(n1061), .ZN(n962) );
  XNOR2_X1 U563 ( .A(n657), .B(n277), .ZN(n724) );
  XNOR2_X1 U564 ( .A(n733), .B(n734), .ZN(n657) );
  NOR2_X1 U565 ( .A1(n386), .A2(n432), .ZN(n389) );
  NAND2_X1 U566 ( .A1(n367), .A2(n366), .ZN(n354) );
  INV_X1 U567 ( .A(n2124), .ZN(n1849) );
  NAND2_X1 U568 ( .A1(n1536), .A2(n1535), .ZN(n1540) );
  OR2_X1 U569 ( .A1(n1538), .A2(n1537), .ZN(n1535) );
  NAND2_X1 U570 ( .A1(n1538), .A2(n1537), .ZN(n1539) );
  XNOR2_X1 U571 ( .A(n1324), .B(fmem_data[31]), .ZN(n1511) );
  XNOR2_X1 U572 ( .A(n1595), .B(n1534), .ZN(n1563) );
  XNOR2_X1 U573 ( .A(n1592), .B(n1593), .ZN(n1534) );
  XNOR2_X1 U574 ( .A(n1324), .B(fmem_data[7]), .ZN(n1236) );
  XNOR2_X1 U575 ( .A(n1324), .B(fmem_data[10]), .ZN(n1192) );
  NAND2_X1 U576 ( .A1(n1628), .A2(n1627), .ZN(n1938) );
  NAND2_X1 U577 ( .A1(n1626), .A2(n1625), .ZN(n1627) );
  OAI21_X1 U578 ( .B1(n1626), .B2(n1625), .A(n1624), .ZN(n1628) );
  NAND2_X1 U579 ( .A1(n1621), .A2(n1620), .ZN(n1622) );
  XNOR2_X1 U580 ( .A(n1334), .B(n200), .ZN(n1152) );
  NAND2_X1 U581 ( .A1(n1553), .A2(n1552), .ZN(n1554) );
  NOR2_X1 U582 ( .A1(n1553), .A2(n1552), .ZN(n1556) );
  INV_X1 U583 ( .A(n1551), .ZN(n1555) );
  INV_X1 U584 ( .A(n1014), .ZN(n1019) );
  NOR2_X1 U585 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  NAND2_X1 U586 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  BUF_X1 U587 ( .A(n1571), .Z(n1547) );
  OR2_X1 U588 ( .A1(n1769), .A2(n1768), .ZN(n1771) );
  AND2_X1 U589 ( .A1(n1910), .A2(n1909), .ZN(n1983) );
  NAND2_X1 U590 ( .A1(n1299), .A2(n1298), .ZN(n1136) );
  AND2_X1 U591 ( .A1(n1948), .A2(n1947), .ZN(n1976) );
  NAND2_X1 U592 ( .A1(n1421), .A2(n1420), .ZN(n1404) );
  NOR2_X1 U593 ( .A1(n1421), .A2(n1420), .ZN(n1405) );
  INV_X1 U594 ( .A(n1422), .ZN(n1406) );
  XNOR2_X1 U595 ( .A(n1431), .B(n1430), .ZN(n1432) );
  OAI21_X1 U596 ( .B1(n1037), .B2(n630), .A(n629), .ZN(n654) );
  XNOR2_X1 U597 ( .A(n446), .B(n445), .ZN(n465) );
  XNOR2_X1 U598 ( .A(n444), .B(n443), .ZN(n446) );
  INV_X1 U599 ( .A(n3697), .ZN(n3896) );
  NOR2_X1 U600 ( .A1(xmem_addr[5]), .A2(n4081), .ZN(n3779) );
  INV_X1 U601 ( .A(n2236), .ZN(n3714) );
  NOR2_X1 U602 ( .A1(xmem_addr[5]), .A2(xmem_addr[4]), .ZN(n3728) );
  INV_X1 U603 ( .A(n2237), .ZN(n3710) );
  OAI21_X1 U604 ( .B1(n1004), .B2(n1003), .A(n1002), .ZN(n1465) );
  NAND2_X1 U605 ( .A1(n1052), .A2(n1051), .ZN(n1086) );
  NAND2_X1 U606 ( .A1(n1048), .A2(n1047), .ZN(n1052) );
  NAND2_X1 U607 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  XNOR2_X1 U608 ( .A(n974), .B(n973), .ZN(n997) );
  XNOR2_X1 U609 ( .A(n972), .B(n971), .ZN(n974) );
  NAND2_X1 U610 ( .A1(n967), .A2(n966), .ZN(n996) );
  NAND2_X1 U611 ( .A1(n965), .A2(n993), .ZN(n967) );
  XNOR2_X1 U612 ( .A(n1064), .B(n1063), .ZN(n1075) );
  NAND2_X1 U613 ( .A1(n735), .A2(n734), .ZN(n736) );
  INV_X1 U614 ( .A(n838), .ZN(n834) );
  INV_X1 U615 ( .A(n837), .ZN(n835) );
  NAND2_X1 U616 ( .A1(n746), .A2(n745), .ZN(n754) );
  NAND2_X1 U617 ( .A1(n742), .A2(n741), .ZN(n746) );
  NAND2_X1 U618 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U619 ( .A(n742), .B(n685), .ZN(n753) );
  NAND3_X1 U620 ( .A1(xmem_addr[3]), .A2(n3728), .A3(n3896), .ZN(n3750) );
  NAND3_X1 U621 ( .A1(xmem_addr[3]), .A2(n3779), .A3(n3896), .ZN(n3801) );
  NAND3_X1 U622 ( .A1(n3779), .A2(n3896), .A3(n4083), .ZN(n3775) );
  NAND2_X1 U623 ( .A1(s_ready_x), .A2(s_valid_x), .ZN(n3697) );
  NAND2_X1 U624 ( .A1(xmem_addr[2]), .A2(n3779), .ZN(n2267) );
  NAND2_X1 U625 ( .A1(n3728), .A2(n4105), .ZN(n2263) );
  BUF_X1 U626 ( .A(n3177), .Z(n3583) );
  BUF_X1 U627 ( .A(n3208), .Z(n3601) );
  BUF_X1 U628 ( .A(n3617), .Z(n3245) );
  BUF_X1 U629 ( .A(n3603), .Z(n3096) );
  BUF_X1 U630 ( .A(n3592), .Z(n3190) );
  BUF_X1 U631 ( .A(n3567), .Z(n3225) );
  XNOR2_X1 U632 ( .A(n1301), .B(n1300), .ZN(n1347) );
  XNOR2_X1 U633 ( .A(n1299), .B(n1298), .ZN(n1300) );
  NAND2_X1 U634 ( .A1(n1468), .A2(n1467), .ZN(n1290) );
  INV_X1 U635 ( .A(n1793), .ZN(n1749) );
  OR2_X1 U636 ( .A1(n1753), .A2(n1752), .ZN(n1599) );
  XNOR2_X1 U637 ( .A(n939), .B(n1048), .ZN(n1085) );
  NAND2_X1 U638 ( .A1(n976), .A2(n975), .ZN(n1084) );
  NAND2_X1 U639 ( .A1(n996), .A2(n995), .ZN(n975) );
  OAI21_X1 U640 ( .B1(n996), .B2(n995), .A(n997), .ZN(n976) );
  NAND2_X1 U641 ( .A1(n987), .A2(n986), .ZN(n1073) );
  NAND2_X1 U642 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U643 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U644 ( .A1(n833), .A2(n836), .ZN(n840) );
  NAND2_X1 U645 ( .A1(n835), .A2(n834), .ZN(n836) );
  OAI21_X1 U646 ( .B1(n389), .B2(n388), .A(n387), .ZN(n700) );
  INV_X1 U647 ( .A(n434), .ZN(n388) );
  NAND2_X1 U648 ( .A1(n386), .A2(n432), .ZN(n387) );
  NOR2_X1 U649 ( .A1(n1827), .A2(reset), .ZN(n3291) );
  NAND2_X1 U650 ( .A1(m_valid_y), .A2(m_ready_y), .ZN(n4009) );
  AND2_X1 U651 ( .A1(n3293), .A2(n3290), .ZN(n3306) );
  BUF_X1 U652 ( .A(n3581), .Z(n3193) );
  BUF_X1 U653 ( .A(n3219), .Z(n3619) );
  BUF_X1 U654 ( .A(n3579), .Z(n3220) );
  CLKBUF_X1 U655 ( .A(n2972), .Z(n3593) );
  NAND2_X1 U656 ( .A1(n1861), .A2(n1860), .ZN(n1863) );
  NAND2_X1 U657 ( .A1(n302), .A2(n1859), .ZN(n1861) );
  INV_X1 U658 ( .A(n2091), .ZN(n3645) );
  OR2_X1 U659 ( .A1(\mac_unit_inst/adder_reg [25]), .A2(
        \mac_unit_inst/x_mult_f_reg [25]), .ZN(n3470) );
  NOR2_X1 U660 ( .A1(n1917), .A2(n1916), .ZN(n308) );
  INV_X2 U661 ( .A(n317), .ZN(n3594) );
  NAND2_X2 U662 ( .A1(n3306), .A2(n3305), .ZN(n3492) );
  NOR2_X1 U663 ( .A1(n1920), .A2(n1919), .ZN(n310) );
  NOR2_X1 U664 ( .A1(n1927), .A2(n1926), .ZN(n311) );
  XOR2_X1 U665 ( .A(n1920), .B(n1919), .Z(n314) );
  INV_X2 U666 ( .A(n3082), .ZN(n3582) );
  XNOR2_X1 U667 ( .A(n4050), .B(n4051), .ZN(n423) );
  AND2_X1 U668 ( .A1(n441), .A2(n442), .ZN(n316) );
  OR2_X1 U669 ( .A1(n2258), .A2(n2261), .ZN(n317) );
  XOR2_X1 U670 ( .A(n1930), .B(n1929), .Z(n332) );
  AND2_X1 U671 ( .A1(n1946), .A2(n1945), .ZN(n334) );
  XOR2_X1 U672 ( .A(n1913), .B(n1912), .Z(n335) );
  AND2_X1 U673 ( .A1(n2028), .A2(n1874), .ZN(n336) );
  XOR2_X1 U674 ( .A(n1917), .B(n1916), .Z(n337) );
  XOR2_X1 U675 ( .A(n1927), .B(n1926), .Z(n338) );
  NOR2_X1 U676 ( .A1(n1915), .A2(n1914), .ZN(n340) );
  OR2_X1 U677 ( .A1(n1485), .A2(n1484), .ZN(n341) );
  OR2_X1 U678 ( .A1(n2223), .A2(n4137), .ZN(n342) );
  OR2_X1 U679 ( .A1(n2223), .A2(n4132), .ZN(n343) );
  OR2_X1 U680 ( .A1(n2223), .A2(n4134), .ZN(n344) );
  OR2_X1 U681 ( .A1(n2223), .A2(n4135), .ZN(n345) );
  OR2_X1 U682 ( .A1(n2223), .A2(n4133), .ZN(n346) );
  XNOR2_X1 U685 ( .A(n886), .B(n228), .ZN(n390) );
  XNOR2_X1 U686 ( .A(n886), .B(fmem_data[4]), .ZN(n408) );
  OAI22_X1 U687 ( .A1(n297), .A2(n390), .B1(n408), .B2(n1010), .ZN(n367) );
  INV_X1 U688 ( .A(n367), .ZN(n350) );
  XOR2_X1 U689 ( .A(xmem_data[8]), .B(xmem_data[9]), .Z(n348) );
  NAND2_X1 U690 ( .A1(n348), .A2(n385), .ZN(n393) );
  BUF_X4 U691 ( .A(xmem_data[9]), .Z(n890) );
  XNOR2_X1 U692 ( .A(fmem_data[5]), .B(n890), .ZN(n394) );
  XNOR2_X1 U693 ( .A(fmem_data[6]), .B(n890), .ZN(n411) );
  OAI22_X1 U694 ( .A1(n931), .A2(n394), .B1(n1036), .B2(n411), .ZN(n366) );
  INV_X1 U695 ( .A(n366), .ZN(n349) );
  NAND2_X1 U696 ( .A1(n350), .A2(n349), .ZN(n353) );
  NAND2_X1 U697 ( .A1(n351), .A2(n352), .ZN(n373) );
  BUF_X4 U698 ( .A(xmem_data[3]), .Z(n709) );
  XNOR2_X1 U699 ( .A(n203), .B(n709), .ZN(n374) );
  OAI22_X1 U700 ( .A1(n711), .A2(n374), .B1(n401), .B2(n774), .ZN(n382) );
  NAND2_X1 U701 ( .A1(xmem_data[1]), .A2(n315), .ZN(n357) );
  BUF_X2 U702 ( .A(n357), .Z(n642) );
  XNOR2_X1 U703 ( .A(fmem_data[12]), .B(n225), .ZN(n384) );
  XNOR2_X1 U704 ( .A(fmem_data[13]), .B(n225), .ZN(n358) );
  OAI22_X1 U705 ( .A1(n642), .A2(n384), .B1(n358), .B2(n315), .ZN(n381) );
  NAND2_X1 U706 ( .A1(n353), .A2(n369), .ZN(n355) );
  NAND2_X1 U707 ( .A1(n355), .A2(n354), .ZN(n660) );
  INV_X1 U708 ( .A(n141), .ZN(n356) );
  AND2_X1 U709 ( .A1(n284), .A2(n356), .ZN(n372) );
  XNOR2_X1 U710 ( .A(fmem_data[14]), .B(n226), .ZN(n410) );
  OAI22_X1 U711 ( .A1(n547), .A2(n358), .B1(n410), .B2(n315), .ZN(n371) );
  XOR2_X1 U712 ( .A(xmem_data[5]), .B(xmem_data[4]), .Z(n359) );
  XNOR2_X1 U713 ( .A(xmem_data[4]), .B(xmem_data[3]), .ZN(n360) );
  NAND2_X1 U714 ( .A1(n359), .A2(n360), .ZN(n383) );
  XNOR2_X1 U715 ( .A(n791), .B(n184), .ZN(n391) );
  XNOR2_X1 U716 ( .A(n791), .B(fmem_data[10]), .ZN(n405) );
  OAI22_X1 U717 ( .A1(n801), .A2(n391), .B1(n405), .B2(n857), .ZN(n370) );
  NAND2_X1 U718 ( .A1(n362), .A2(n361), .ZN(n402) );
  XNOR2_X1 U719 ( .A(fmem_data[2]), .B(n252), .ZN(n403) );
  XNOR2_X1 U720 ( .A(xmem_data[11]), .B(xmem_data[12]), .ZN(n375) );
  XNOR2_X1 U721 ( .A(n229), .B(n252), .ZN(n632) );
  OAI22_X1 U722 ( .A1(n1246), .A2(n403), .B1(n1233), .B2(n632), .ZN(n666) );
  XNOR2_X1 U723 ( .A(n4055), .B(n4067), .ZN(n378) );
  NAND2_X1 U724 ( .A1(n378), .A2(n363), .ZN(n377) );
  BUF_X2 U725 ( .A(n377), .Z(n875) );
  XNOR2_X1 U726 ( .A(fmem_data[8]), .B(n849), .ZN(n399) );
  XNOR2_X1 U727 ( .A(fmem_data[9]), .B(n849), .ZN(n636) );
  OAI22_X1 U728 ( .A1(n875), .A2(n399), .B1(n871), .B2(n636), .ZN(n665) );
  NAND2_X1 U729 ( .A1(n406), .A2(n364), .ZN(n723) );
  XNOR2_X1 U730 ( .A(n284), .B(n1269), .ZN(n365) );
  XNOR2_X1 U731 ( .A(fmem_data[1]), .B(n1269), .ZN(n637) );
  OAI22_X1 U732 ( .A1(n723), .A2(n365), .B1(n141), .B2(n637), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U734 ( .A(n369), .B(n368), .ZN(n433) );
  FA_X1 U735 ( .A(n372), .B(n371), .CI(n370), .CO(n659), .S(n432) );
  XNOR2_X1 U736 ( .A(fmem_data[9]), .B(n709), .ZN(n421) );
  OAI22_X1 U737 ( .A1(n138), .A2(n421), .B1(n374), .B2(n774), .ZN(n444) );
  INV_X1 U738 ( .A(n1249), .ZN(n376) );
  AND2_X1 U739 ( .A1(n286), .A2(n376), .ZN(n443) );
  BUF_X2 U740 ( .A(n377), .Z(n870) );
  XNOR2_X1 U741 ( .A(fmem_data[5]), .B(n279), .ZN(n427) );
  XNOR2_X1 U742 ( .A(fmem_data[6]), .B(n279), .ZN(n397) );
  OAI22_X1 U743 ( .A1(n870), .A2(n427), .B1(n871), .B2(n397), .ZN(n445) );
  OAI21_X1 U744 ( .B1(n444), .B2(n443), .A(n445), .ZN(n380) );
  NAND2_X1 U745 ( .A1(n444), .A2(n443), .ZN(n379) );
  NAND2_X1 U746 ( .A1(n380), .A2(n379), .ZN(n438) );
  HA_X1 U747 ( .A(n382), .B(n381), .CO(n369), .S(n437) );
  XNOR2_X1 U748 ( .A(n261), .B(n238), .ZN(n440) );
  XNOR2_X1 U749 ( .A(n791), .B(fmem_data[8]), .ZN(n392) );
  OAI22_X1 U750 ( .A1(n858), .A2(n440), .B1(n392), .B2(n857), .ZN(n449) );
  XNOR2_X1 U751 ( .A(fmem_data[11]), .B(n639), .ZN(n422) );
  OAI22_X1 U752 ( .A1(n547), .A2(n422), .B1(n384), .B2(n315), .ZN(n448) );
  XNOR2_X1 U753 ( .A(n229), .B(n189), .ZN(n439) );
  XNOR2_X1 U754 ( .A(fmem_data[4]), .B(n890), .ZN(n395) );
  OAI22_X1 U755 ( .A1(n1037), .A2(n439), .B1(n929), .B2(n395), .ZN(n447) );
  BUF_X2 U756 ( .A(xmem_data[11]), .Z(n1231) );
  XNOR2_X1 U757 ( .A(n1231), .B(fmem_data[2]), .ZN(n424) );
  OAI22_X1 U758 ( .A1(n296), .A2(n424), .B1(n390), .B2(n1010), .ZN(n417) );
  OAI22_X1 U759 ( .A1(n858), .A2(n392), .B1(n391), .B2(n857), .ZN(n416) );
  OAI22_X1 U760 ( .A1(n1037), .A2(n395), .B1(n1036), .B2(n394), .ZN(n415) );
  XNOR2_X1 U761 ( .A(n287), .B(n252), .ZN(n396) );
  XNOR2_X1 U762 ( .A(fmem_data[1]), .B(n252), .ZN(n404) );
  OAI22_X1 U763 ( .A1(n1246), .A2(n396), .B1(n1249), .B2(n404), .ZN(n420) );
  XNOR2_X1 U764 ( .A(fmem_data[7]), .B(n279), .ZN(n400) );
  OAI22_X1 U765 ( .A1(n870), .A2(n397), .B1(n871), .B2(n400), .ZN(n419) );
  OR2_X1 U766 ( .A1(n285), .A2(n214), .ZN(n398) );
  OAI22_X1 U767 ( .A1(n1246), .A2(n214), .B1(n1249), .B2(n398), .ZN(n418) );
  OAI22_X1 U768 ( .A1(n875), .A2(n400), .B1(n871), .B2(n399), .ZN(n414) );
  OAI22_X1 U769 ( .A1(n711), .A2(n401), .B1(n409), .B2(n774), .ZN(n413) );
  BUF_X2 U770 ( .A(n402), .Z(n1246) );
  OAI22_X1 U771 ( .A1(n1246), .A2(n404), .B1(n1249), .B2(n403), .ZN(n412) );
  XNOR2_X1 U772 ( .A(n791), .B(fmem_data[11]), .ZN(n638) );
  OAI22_X1 U773 ( .A1(n801), .A2(n405), .B1(n638), .B2(n857), .ZN(n671) );
  OR2_X1 U774 ( .A1(n286), .A2(n4053), .ZN(n407) );
  OAI22_X1 U775 ( .A1(n201), .A2(n4053), .B1(n219), .B2(n407), .ZN(n670) );
  XNOR2_X1 U776 ( .A(n1231), .B(fmem_data[5]), .ZN(n631) );
  OAI22_X1 U777 ( .A1(n296), .A2(n408), .B1(n631), .B2(n1010), .ZN(n669) );
  XNOR2_X1 U778 ( .A(fmem_data[13]), .B(n709), .ZN(n634) );
  OAI22_X1 U779 ( .A1(n711), .A2(n409), .B1(n634), .B2(n774), .ZN(n668) );
  XNOR2_X1 U780 ( .A(fmem_data[15]), .B(n225), .ZN(n640) );
  OAI22_X1 U781 ( .A1(n547), .A2(n410), .B1(n640), .B2(n315), .ZN(n667) );
  XNOR2_X1 U782 ( .A(n238), .B(n890), .ZN(n630) );
  OAI22_X1 U783 ( .A1(n1037), .A2(n411), .B1(n1036), .B2(n630), .ZN(n662) );
  FA_X1 U784 ( .A(n414), .B(n413), .CI(n412), .CO(n661), .S(n429) );
  FA_X1 U785 ( .A(n417), .B(n416), .CI(n415), .CO(n431), .S(n452) );
  FA_X1 U786 ( .A(n420), .B(n419), .CI(n418), .CO(n430), .S(n451) );
  XNOR2_X1 U787 ( .A(fmem_data[8]), .B(n709), .ZN(n460) );
  OAI22_X1 U788 ( .A1(n138), .A2(n460), .B1(n421), .B2(n774), .ZN(n442) );
  XNOR2_X1 U789 ( .A(fmem_data[10]), .B(n639), .ZN(n458) );
  OAI22_X1 U790 ( .A1(n642), .A2(n458), .B1(n422), .B2(n315), .ZN(n441) );
  XNOR2_X1 U791 ( .A(n1231), .B(fmem_data[1]), .ZN(n425) );
  OAI22_X1 U792 ( .A1(n296), .A2(n425), .B1(n424), .B2(n1010), .ZN(n454) );
  XNOR2_X1 U793 ( .A(n886), .B(n286), .ZN(n426) );
  OAI22_X1 U794 ( .A1(n296), .A2(n426), .B1(n425), .B2(n1010), .ZN(n463) );
  XNOR2_X1 U795 ( .A(fmem_data[4]), .B(n279), .ZN(n456) );
  OAI22_X1 U796 ( .A1(n870), .A2(n456), .B1(n871), .B2(n427), .ZN(n462) );
  OR2_X1 U797 ( .A1(n284), .A2(n4058), .ZN(n428) );
  OAI22_X1 U798 ( .A1(n297), .A2(n4058), .B1(n428), .B2(n1010), .ZN(n461) );
  FA_X1 U799 ( .A(n431), .B(n430), .CI(n429), .CO(n688), .S(n468) );
  XNOR2_X1 U800 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X1 U801 ( .A(n435), .B(n434), .ZN(n467) );
  FA_X1 U802 ( .A(n438), .B(n437), .CI(n436), .CO(n434), .S(n472) );
  XNOR2_X1 U803 ( .A(fmem_data[2]), .B(n189), .ZN(n457) );
  OAI22_X1 U804 ( .A1(n1037), .A2(n457), .B1(n929), .B2(n439), .ZN(n597) );
  XNOR2_X1 U805 ( .A(n261), .B(fmem_data[6]), .ZN(n455) );
  OAI22_X1 U806 ( .A1(n801), .A2(n455), .B1(n440), .B2(n857), .ZN(n596) );
  XOR2_X1 U807 ( .A(n442), .B(n441), .Z(n595) );
  FA_X1 U808 ( .A(n449), .B(n448), .CI(n447), .CO(n436), .S(n464) );
  FA_X1 U809 ( .A(n452), .B(n451), .CI(n450), .CO(n469), .S(n470) );
  FA_X1 U810 ( .A(n316), .B(n454), .CI(n453), .CO(n450), .S(n606) );
  XNOR2_X1 U811 ( .A(n261), .B(n183), .ZN(n484) );
  OAI22_X1 U812 ( .A1(n858), .A2(n484), .B1(n455), .B2(n857), .ZN(n483) );
  XNOR2_X1 U813 ( .A(n228), .B(n279), .ZN(n485) );
  OAI22_X1 U814 ( .A1(n870), .A2(n485), .B1(n871), .B2(n456), .ZN(n482) );
  XNOR2_X1 U815 ( .A(fmem_data[1]), .B(n890), .ZN(n487) );
  OAI22_X1 U816 ( .A1(n1037), .A2(n487), .B1(n1036), .B2(n457), .ZN(n481) );
  XNOR2_X1 U817 ( .A(fmem_data[9]), .B(n226), .ZN(n477) );
  OAI22_X1 U818 ( .A1(n642), .A2(n477), .B1(n458), .B2(n315), .ZN(n493) );
  INV_X1 U819 ( .A(n1010), .ZN(n459) );
  AND2_X1 U820 ( .A1(n284), .A2(n459), .ZN(n492) );
  XNOR2_X1 U821 ( .A(fmem_data[7]), .B(n709), .ZN(n476) );
  OAI22_X1 U822 ( .A1(n138), .A2(n476), .B1(n460), .B2(n774), .ZN(n491) );
  FA_X1 U823 ( .A(n466), .B(n465), .CI(n464), .CO(n471), .S(n604) );
  NOR2_X1 U824 ( .A1(n620), .A2(n619), .ZN(n1828) );
  INV_X1 U825 ( .A(n1828), .ZN(n3646) );
  FA_X1 U826 ( .A(n467), .B(n468), .CI(n469), .CO(n623), .S(n622) );
  INV_X1 U827 ( .A(n622), .ZN(n474) );
  FA_X1 U828 ( .A(n472), .B(n471), .CI(n470), .CO(n621), .S(n620) );
  INV_X1 U829 ( .A(n621), .ZN(n473) );
  NAND2_X1 U830 ( .A1(n474), .A2(n473), .ZN(n2093) );
  NAND2_X1 U831 ( .A1(n3646), .A2(n2093), .ZN(n475) );
  NOR2_X1 U832 ( .A1(n237), .A2(n475), .ZN(n628) );
  XNOR2_X1 U833 ( .A(fmem_data[6]), .B(n709), .ZN(n480) );
  OAI22_X1 U834 ( .A1(n138), .A2(n480), .B1(n476), .B2(n774), .ZN(n490) );
  XNOR2_X1 U835 ( .A(n258), .B(n226), .ZN(n498) );
  OAI22_X1 U836 ( .A1(n547), .A2(n498), .B1(n477), .B2(n315), .ZN(n489) );
  OR2_X1 U837 ( .A1(n287), .A2(n190), .ZN(n478) );
  OAI22_X1 U838 ( .A1(n1037), .A2(n190), .B1(n929), .B2(n478), .ZN(n502) );
  INV_X1 U839 ( .A(n929), .ZN(n479) );
  AND2_X1 U840 ( .A1(n284), .A2(n479), .ZN(n509) );
  XNOR2_X1 U841 ( .A(fmem_data[5]), .B(n709), .ZN(n499) );
  OAI22_X1 U842 ( .A1(n138), .A2(n499), .B1(n480), .B2(n774), .ZN(n508) );
  XNOR2_X1 U843 ( .A(fmem_data[1]), .B(n279), .ZN(n511) );
  XNOR2_X1 U844 ( .A(fmem_data[2]), .B(n279), .ZN(n486) );
  OAI22_X1 U845 ( .A1(n870), .A2(n511), .B1(n871), .B2(n486), .ZN(n507) );
  FA_X1 U846 ( .A(n483), .B(n482), .CI(n481), .CO(n600), .S(n602) );
  XNOR2_X1 U847 ( .A(n261), .B(fmem_data[4]), .ZN(n497) );
  OAI22_X1 U848 ( .A1(n801), .A2(n497), .B1(n484), .B2(n857), .ZN(n496) );
  OAI22_X1 U849 ( .A1(n870), .A2(n486), .B1(n871), .B2(n485), .ZN(n495) );
  XNOR2_X1 U850 ( .A(n286), .B(n189), .ZN(n488) );
  OAI22_X1 U851 ( .A1(n1037), .A2(n488), .B1(n929), .B2(n487), .ZN(n494) );
  HA_X1 U852 ( .A(n490), .B(n489), .CO(n593), .S(n503) );
  FA_X1 U853 ( .A(n493), .B(n492), .CI(n491), .CO(n599), .S(n592) );
  FA_X1 U854 ( .A(n496), .B(n495), .CI(n494), .CO(n594), .S(n506) );
  XNOR2_X1 U855 ( .A(n261), .B(n228), .ZN(n513) );
  OAI22_X1 U856 ( .A1(n801), .A2(n513), .B1(n497), .B2(n857), .ZN(n516) );
  XNOR2_X1 U857 ( .A(n238), .B(n226), .ZN(n500) );
  OAI22_X1 U858 ( .A1(n642), .A2(n500), .B1(n498), .B2(n315), .ZN(n515) );
  XNOR2_X1 U859 ( .A(n233), .B(n709), .ZN(n518) );
  OAI22_X1 U860 ( .A1(n711), .A2(n518), .B1(n499), .B2(n774), .ZN(n566) );
  XNOR2_X1 U861 ( .A(fmem_data[6]), .B(n226), .ZN(n520) );
  OAI22_X1 U862 ( .A1(n547), .A2(n520), .B1(n500), .B2(n315), .ZN(n565) );
  FA_X1 U863 ( .A(n503), .B(n502), .CI(n501), .CO(n603), .S(n504) );
  FA_X1 U864 ( .A(n506), .B(n505), .CI(n504), .CO(n588), .S(n587) );
  FA_X1 U865 ( .A(n509), .B(n508), .CI(n507), .CO(n501), .S(n579) );
  OR2_X1 U866 ( .A1(n285), .A2(n4068), .ZN(n510) );
  OAI22_X1 U867 ( .A1(n870), .A2(n4068), .B1(n871), .B2(n510), .ZN(n569) );
  XNOR2_X1 U868 ( .A(n287), .B(n279), .ZN(n512) );
  OAI22_X1 U869 ( .A1(n870), .A2(n512), .B1(n871), .B2(n511), .ZN(n568) );
  XNOR2_X1 U870 ( .A(n261), .B(fmem_data[2]), .ZN(n517) );
  OAI22_X1 U871 ( .A1(n858), .A2(n517), .B1(n513), .B2(n857), .ZN(n567) );
  FA_X1 U872 ( .A(n516), .B(n515), .CI(n514), .CO(n505), .S(n577) );
  NOR2_X1 U873 ( .A1(n2179), .A2(n2164), .ZN(n591) );
  XNOR2_X1 U874 ( .A(fmem_data[2]), .B(n709), .ZN(n533) );
  XNOR2_X1 U875 ( .A(n229), .B(n709), .ZN(n519) );
  OAI22_X1 U876 ( .A1(n138), .A2(n533), .B1(n519), .B2(n774), .ZN(n527) );
  XNOR2_X1 U877 ( .A(n233), .B(n225), .ZN(n531) );
  XNOR2_X1 U878 ( .A(n183), .B(n225), .ZN(n521) );
  OAI22_X1 U879 ( .A1(n547), .A2(n531), .B1(n521), .B2(n315), .ZN(n526) );
  XNOR2_X1 U880 ( .A(n261), .B(fmem_data[1]), .ZN(n524) );
  OAI22_X1 U881 ( .A1(n858), .A2(n524), .B1(n517), .B2(n857), .ZN(n571) );
  OAI22_X1 U882 ( .A1(n138), .A2(n519), .B1(n518), .B2(n774), .ZN(n564) );
  OAI22_X1 U883 ( .A1(n642), .A2(n521), .B1(n520), .B2(n315), .ZN(n563) );
  INV_X1 U884 ( .A(n871), .ZN(n522) );
  AND2_X1 U885 ( .A1(n286), .A2(n522), .ZN(n562) );
  OR2_X1 U886 ( .A1(n284), .A2(n4055), .ZN(n523) );
  OAI22_X1 U887 ( .A1(n858), .A2(n4055), .B1(n523), .B2(n857), .ZN(n530) );
  XNOR2_X1 U888 ( .A(n261), .B(n287), .ZN(n525) );
  OAI22_X1 U889 ( .A1(n858), .A2(n525), .B1(n524), .B2(n857), .ZN(n529) );
  HA_X1 U890 ( .A(n527), .B(n526), .CO(n572), .S(n528) );
  NOR2_X1 U891 ( .A1(n560), .A2(n559), .ZN(n1830) );
  FA_X1 U892 ( .A(n530), .B(n529), .CI(n528), .CO(n559), .S(n556) );
  XNOR2_X1 U893 ( .A(n229), .B(n226), .ZN(n539) );
  OAI22_X1 U894 ( .A1(n547), .A2(n539), .B1(n531), .B2(n315), .ZN(n536) );
  INV_X1 U895 ( .A(n857), .ZN(n532) );
  AND2_X1 U896 ( .A1(n284), .A2(n532), .ZN(n535) );
  XNOR2_X1 U897 ( .A(fmem_data[1]), .B(n709), .ZN(n537) );
  OAI22_X1 U898 ( .A1(n138), .A2(n537), .B1(n533), .B2(n774), .ZN(n534) );
  NOR2_X1 U899 ( .A1(n556), .A2(n555), .ZN(n1834) );
  INV_X1 U900 ( .A(n1834), .ZN(n2220) );
  FA_X1 U901 ( .A(n536), .B(n535), .CI(n534), .CO(n555), .S(n554) );
  XNOR2_X1 U902 ( .A(n285), .B(n709), .ZN(n538) );
  OAI22_X1 U903 ( .A1(n138), .A2(n538), .B1(n537), .B2(n774), .ZN(n541) );
  XNOR2_X1 U904 ( .A(fmem_data[2]), .B(n225), .ZN(n543) );
  OAI22_X1 U905 ( .A1(n547), .A2(n543), .B1(n539), .B2(n315), .ZN(n540) );
  NOR2_X1 U906 ( .A1(n554), .A2(n553), .ZN(n1831) );
  HA_X1 U907 ( .A(n541), .B(n540), .CO(n553), .S(n551) );
  OR2_X1 U908 ( .A1(n285), .A2(n198), .ZN(n542) );
  OAI22_X1 U909 ( .A1(n138), .A2(n198), .B1(n542), .B2(n774), .ZN(n550) );
  OR2_X1 U910 ( .A1(n551), .A2(n550), .ZN(n2213) );
  XNOR2_X1 U911 ( .A(fmem_data[1]), .B(n225), .ZN(n546) );
  OAI22_X1 U912 ( .A1(n642), .A2(n546), .B1(n543), .B2(n315), .ZN(n549) );
  INV_X1 U913 ( .A(n774), .ZN(n544) );
  AND2_X1 U914 ( .A1(n287), .A2(n544), .ZN(n548) );
  NOR2_X1 U915 ( .A1(n549), .A2(n548), .ZN(n2204) );
  OR2_X1 U916 ( .A1(n286), .A2(n339), .ZN(n545) );
  NAND2_X1 U917 ( .A1(n545), .A2(n547), .ZN(n2191) );
  OAI22_X1 U918 ( .A1(n547), .A2(n286), .B1(n546), .B2(n315), .ZN(n2190) );
  NAND2_X1 U919 ( .A1(n2191), .A2(n2190), .ZN(n2207) );
  NAND2_X1 U920 ( .A1(n549), .A2(n548), .ZN(n2205) );
  OAI21_X1 U921 ( .B1(n2204), .B2(n2207), .A(n2205), .ZN(n2214) );
  NAND2_X1 U922 ( .A1(n551), .A2(n550), .ZN(n2212) );
  INV_X1 U923 ( .A(n2212), .ZN(n552) );
  AOI21_X1 U924 ( .B1(n2213), .B2(n2214), .A(n552), .ZN(n1832) );
  NAND2_X1 U925 ( .A1(n554), .A2(n553), .ZN(n2196) );
  OAI21_X1 U926 ( .B1(n1831), .B2(n1832), .A(n2196), .ZN(n558) );
  NAND2_X1 U927 ( .A1(n556), .A2(n555), .ZN(n2219) );
  INV_X1 U928 ( .A(n2219), .ZN(n557) );
  AOI21_X1 U929 ( .B1(n2220), .B2(n558), .A(n557), .ZN(n561) );
  NAND2_X1 U930 ( .A1(n560), .A2(n559), .ZN(n2113) );
  OAI21_X1 U931 ( .B1(n1830), .B2(n561), .A(n2113), .ZN(n576) );
  FA_X1 U932 ( .A(n564), .B(n563), .CI(n562), .CO(n582), .S(n570) );
  HA_X1 U933 ( .A(n566), .B(n565), .CO(n514), .S(n581) );
  FA_X1 U934 ( .A(n569), .B(n568), .CI(n567), .CO(n578), .S(n580) );
  FA_X1 U935 ( .A(n572), .B(n571), .CI(n570), .CO(n573), .S(n560) );
  NOR2_X1 U936 ( .A1(n574), .A2(n573), .ZN(n1836) );
  INV_X1 U937 ( .A(n1836), .ZN(n2107) );
  NAND2_X1 U938 ( .A1(n574), .A2(n573), .ZN(n2106) );
  INV_X1 U939 ( .A(n2106), .ZN(n575) );
  AOI21_X1 U940 ( .B1(n576), .B2(n2107), .A(n575), .ZN(n585) );
  FA_X1 U941 ( .A(n579), .B(n578), .CI(n577), .CO(n586), .S(n584) );
  FA_X1 U942 ( .A(n582), .B(n581), .CI(n580), .CO(n583), .S(n574) );
  NOR2_X1 U943 ( .A1(n584), .A2(n583), .ZN(n3651) );
  NAND2_X1 U944 ( .A1(n584), .A2(n583), .ZN(n3652) );
  OAI21_X1 U945 ( .B1(n585), .B2(n3651), .A(n3652), .ZN(n2168) );
  NAND2_X1 U946 ( .A1(n587), .A2(n586), .ZN(n2165) );
  NAND2_X1 U947 ( .A1(n589), .A2(n588), .ZN(n2180) );
  OAI21_X1 U948 ( .B1(n2179), .B2(n2165), .A(n2180), .ZN(n590) );
  AOI21_X1 U949 ( .B1(n591), .B2(n2168), .A(n590), .ZN(n618) );
  FA_X1 U950 ( .A(n594), .B(n593), .CI(n592), .CO(n609), .S(n601) );
  FA_X1 U951 ( .A(n597), .B(n596), .CI(n595), .CO(n466), .S(n608) );
  FA_X1 U952 ( .A(n600), .B(n599), .CI(n598), .CO(n605), .S(n607) );
  FA_X1 U953 ( .A(n603), .B(n602), .CI(n601), .CO(n610), .S(n589) );
  NOR2_X1 U954 ( .A1(n611), .A2(n610), .ZN(n2082) );
  INV_X1 U955 ( .A(n2082), .ZN(n2100) );
  FA_X1 U956 ( .A(n606), .B(n605), .CI(n604), .CO(n619), .S(n613) );
  FA_X1 U957 ( .A(n609), .B(n608), .CI(n607), .CO(n612), .S(n611) );
  OR2_X2 U958 ( .A1(n613), .A2(n612), .ZN(n2084) );
  NAND2_X1 U959 ( .A1(n2100), .A2(n2084), .ZN(n617) );
  NAND2_X1 U960 ( .A1(n611), .A2(n610), .ZN(n2099) );
  INV_X1 U961 ( .A(n2099), .ZN(n615) );
  NAND2_X1 U962 ( .A1(n613), .A2(n612), .ZN(n2083) );
  INV_X1 U963 ( .A(n2083), .ZN(n614) );
  AOI21_X1 U964 ( .B1(n2084), .B2(n615), .A(n614), .ZN(n616) );
  OAI21_X1 U965 ( .B1(n618), .B2(n617), .A(n616), .ZN(n627) );
  AND2_X1 U966 ( .A1(n620), .A2(n619), .ZN(n2091) );
  AOI21_X1 U967 ( .B1(n2093), .B2(n2091), .A(n181), .ZN(n625) );
  NAND2_X1 U968 ( .A1(n624), .A2(n623), .ZN(n2157) );
  OAI21_X1 U969 ( .B1(n625), .B2(n1829), .A(n2157), .ZN(n626) );
  AOI21_X1 U970 ( .B1(n627), .B2(n628), .A(n626), .ZN(n760) );
  XNOR2_X1 U971 ( .A(fmem_data[8]), .B(n890), .ZN(n680) );
  OR2_X1 U972 ( .A1(n929), .A2(n680), .ZN(n629) );
  XNOR2_X1 U973 ( .A(n1231), .B(fmem_data[6]), .ZN(n677) );
  OAI22_X1 U974 ( .A1(n296), .A2(n631), .B1(n677), .B2(n1010), .ZN(n652) );
  XNOR2_X1 U975 ( .A(fmem_data[4]), .B(n252), .ZN(n678) );
  OAI22_X1 U976 ( .A1(n1246), .A2(n632), .B1(n1249), .B2(n678), .ZN(n653) );
  XNOR2_X1 U977 ( .A(n652), .B(n653), .ZN(n633) );
  XNOR2_X1 U978 ( .A(n633), .B(n654), .ZN(n691) );
  XNOR2_X1 U979 ( .A(fmem_data[14]), .B(n709), .ZN(n646) );
  OAI22_X1 U980 ( .A1(n711), .A2(n634), .B1(n646), .B2(n774), .ZN(n651) );
  INV_X1 U981 ( .A(n1353), .ZN(n635) );
  AND2_X1 U982 ( .A1(n284), .A2(n635), .ZN(n650) );
  XNOR2_X1 U983 ( .A(fmem_data[10]), .B(n849), .ZN(n645) );
  OAI22_X1 U984 ( .A1(n870), .A2(n636), .B1(n871), .B2(n645), .ZN(n649) );
  XNOR2_X1 U985 ( .A(fmem_data[2]), .B(n1113), .ZN(n679) );
  OAI22_X1 U986 ( .A1(n201), .A2(n637), .B1(n141), .B2(n679), .ZN(n648) );
  XNOR2_X1 U987 ( .A(n791), .B(fmem_data[12]), .ZN(n644) );
  OAI22_X1 U988 ( .A1(n858), .A2(n638), .B1(n644), .B2(n857), .ZN(n647) );
  XNOR2_X1 U989 ( .A(fmem_data[31]), .B(n226), .ZN(n641) );
  AOI21_X1 U990 ( .B1(n642), .B2(n315), .A(n641), .ZN(n643) );
  INV_X1 U991 ( .A(n643), .ZN(n732) );
  XNOR2_X1 U992 ( .A(n261), .B(n194), .ZN(n729) );
  OAI22_X1 U993 ( .A1(n858), .A2(n644), .B1(n729), .B2(n857), .ZN(n731) );
  XNOR2_X1 U994 ( .A(fmem_data[11]), .B(n279), .ZN(n712) );
  OAI22_X1 U995 ( .A1(n870), .A2(n645), .B1(n871), .B2(n712), .ZN(n708) );
  XNOR2_X1 U996 ( .A(fmem_data[15]), .B(n709), .ZN(n710) );
  OAI22_X1 U997 ( .A1(n138), .A2(n646), .B1(n710), .B2(n774), .ZN(n707) );
  XNOR2_X1 U998 ( .A(n708), .B(n707), .ZN(n730) );
  OAI21_X1 U999 ( .B1(n653), .B2(n654), .A(n652), .ZN(n656) );
  NAND2_X1 U1000 ( .A1(n656), .A2(n655), .ZN(n735) );
  FA_X1 U1001 ( .A(n660), .B(n659), .CI(n658), .CO(n694), .S(n701) );
  FA_X1 U1002 ( .A(n663), .B(n662), .CI(n661), .CO(n692), .S(n686) );
  FA_X1 U1003 ( .A(n664), .B(n665), .CI(n666), .CO(n676), .S(n658) );
  HA_X1 U1004 ( .A(n668), .B(n667), .CO(n675), .S(n663) );
  FA_X1 U1005 ( .A(n671), .B(n670), .CI(n669), .CO(n674), .S(n687) );
  OAI21_X1 U1006 ( .B1(n694), .B2(n692), .A(n693), .ZN(n673) );
  NAND2_X1 U1007 ( .A1(n694), .A2(n692), .ZN(n672) );
  NAND2_X1 U1008 ( .A1(n673), .A2(n672), .ZN(n744) );
  FA_X1 U1009 ( .A(n676), .B(n675), .CI(n674), .CO(n705), .S(n693) );
  XNOR2_X1 U1010 ( .A(n886), .B(fmem_data[7]), .ZN(n720) );
  OAI22_X1 U1011 ( .A1(n297), .A2(n677), .B1(n720), .B2(n1010), .ZN(n719) );
  XNOR2_X1 U1012 ( .A(fmem_data[5]), .B(n252), .ZN(n721) );
  OAI22_X1 U1013 ( .A1(n1246), .A2(n678), .B1(n1233), .B2(n721), .ZN(n718) );
  XNOR2_X1 U1014 ( .A(n228), .B(n1113), .ZN(n722) );
  OAI22_X1 U1015 ( .A1(n723), .A2(n679), .B1(n141), .B2(n722), .ZN(n717) );
  XNOR2_X1 U1016 ( .A(fmem_data[9]), .B(n890), .ZN(n727) );
  OAI22_X1 U1017 ( .A1(n931), .A2(n680), .B1(n1036), .B2(n727), .ZN(n716) );
  NAND2_X1 U1018 ( .A1(n681), .A2(n788), .ZN(n925) );
  BUF_X2 U1019 ( .A(n925), .Z(n1356) );
  BUF_X4 U1020 ( .A(xmem_data[17]), .Z(n1266) );
  OR2_X1 U1021 ( .A1(n285), .A2(n180), .ZN(n682) );
  OAI22_X1 U1022 ( .A1(n1356), .A2(n180), .B1(n682), .B2(n1353), .ZN(n715) );
  XNOR2_X1 U1023 ( .A(n1266), .B(n286), .ZN(n683) );
  XNOR2_X1 U1024 ( .A(n1266), .B(fmem_data[1]), .ZN(n728) );
  OAI22_X1 U1025 ( .A1(n1356), .A2(n683), .B1(n728), .B2(n1353), .ZN(n714) );
  XNOR2_X1 U1026 ( .A(n744), .B(n743), .ZN(n685) );
  FA_X1 U1027 ( .A(n688), .B(n687), .CI(n686), .CO(n698), .S(n699) );
  FA_X1 U1028 ( .A(n691), .B(n690), .CI(n689), .CO(n726), .S(n697) );
  XNOR2_X1 U1029 ( .A(n693), .B(n692), .ZN(n695) );
  XNOR2_X1 U1030 ( .A(n695), .B(n694), .ZN(n696) );
  FA_X1 U1031 ( .A(n698), .B(n697), .CI(n696), .CO(n752), .S(n751) );
  FA_X1 U1032 ( .A(n701), .B(n700), .CI(n699), .CO(n750), .S(n624) );
  NOR2_X1 U1033 ( .A1(n751), .A2(n750), .ZN(n2139) );
  NOR2_X1 U1034 ( .A1(n1846), .A2(n2139), .ZN(n749) );
  OR2_X1 U1035 ( .A1(n703), .A2(n702), .ZN(n704) );
  AOI22_X1 U1036 ( .A1(n705), .A2(n704), .B1(n703), .B2(n702), .ZN(n706) );
  INV_X1 U1037 ( .A(n706), .ZN(n823) );
  OR2_X1 U1038 ( .A1(n708), .A2(n707), .ZN(n816) );
  XNOR2_X1 U1039 ( .A(fmem_data[31]), .B(n709), .ZN(n773) );
  OAI22_X1 U1040 ( .A1(n773), .A2(n774), .B1(n138), .B2(n710), .ZN(n815) );
  XNOR2_X1 U1041 ( .A(fmem_data[12]), .B(n279), .ZN(n762) );
  OAI22_X1 U1042 ( .A1(n870), .A2(n712), .B1(n871), .B2(n762), .ZN(n777) );
  XNOR2_X1 U1043 ( .A(n4059), .B(n4060), .ZN(n764) );
  INV_X1 U1044 ( .A(n1253), .ZN(n713) );
  AND2_X1 U1045 ( .A1(n286), .A2(n713), .ZN(n776) );
  XNOR2_X1 U1046 ( .A(n777), .B(n776), .ZN(n814) );
  FA_X1 U1047 ( .A(n716), .B(n715), .CI(n714), .CO(n819), .S(n702) );
  FA_X1 U1048 ( .A(n719), .B(n718), .CI(n717), .CO(n818), .S(n703) );
  XNOR2_X1 U1049 ( .A(n886), .B(fmem_data[8]), .ZN(n770) );
  OAI22_X1 U1050 ( .A1(n295), .A2(n720), .B1(n770), .B2(n1010), .ZN(n780) );
  XNOR2_X1 U1051 ( .A(fmem_data[6]), .B(n1245), .ZN(n761) );
  OAI22_X1 U1052 ( .A1(n721), .A2(n1251), .B1(n1249), .B2(n761), .ZN(n779) );
  XNOR2_X1 U1053 ( .A(fmem_data[4]), .B(n1113), .ZN(n772) );
  OAI22_X1 U1054 ( .A1(n201), .A2(n722), .B1(n219), .B2(n772), .ZN(n778) );
  FA_X1 U1055 ( .A(n726), .B(n725), .CI(n724), .CO(n838), .S(n742) );
  XNOR2_X1 U1056 ( .A(fmem_data[10]), .B(n890), .ZN(n796) );
  OAI22_X1 U1057 ( .A1(n1037), .A2(n727), .B1(n929), .B2(n796), .ZN(n769) );
  XNOR2_X1 U1058 ( .A(n1266), .B(fmem_data[2]), .ZN(n798) );
  OAI22_X1 U1059 ( .A1(n1356), .A2(n728), .B1(n798), .B2(n1353), .ZN(n768) );
  XNOR2_X1 U1060 ( .A(n261), .B(fmem_data[14]), .ZN(n800) );
  OAI22_X1 U1061 ( .A1(n801), .A2(n729), .B1(n800), .B2(n857), .ZN(n767) );
  FA_X1 U1062 ( .A(n732), .B(n731), .CI(n730), .CO(n782), .S(n725) );
  OAI21_X1 U1063 ( .B1(n735), .B2(n734), .A(n733), .ZN(n737) );
  NAND2_X1 U1064 ( .A1(n737), .A2(n736), .ZN(n781) );
  XNOR2_X1 U1065 ( .A(n838), .B(n837), .ZN(n738) );
  XNOR2_X1 U1066 ( .A(n738), .B(n833), .ZN(n755) );
  INV_X1 U1067 ( .A(n755), .ZN(n748) );
  INV_X1 U1068 ( .A(n744), .ZN(n739) );
  NAND2_X1 U1069 ( .A1(n744), .A2(n743), .ZN(n745) );
  INV_X1 U1070 ( .A(n754), .ZN(n747) );
  NAND2_X1 U1071 ( .A1(n749), .A2(n2124), .ZN(n759) );
  NAND2_X1 U1072 ( .A1(n751), .A2(n750), .ZN(n3640) );
  NAND2_X1 U1073 ( .A1(n753), .A2(n752), .ZN(n2140) );
  OAI21_X1 U1074 ( .B1(n1846), .B2(n3640), .A(n2140), .ZN(n757) );
  NAND2_X1 U1075 ( .A1(n755), .A2(n754), .ZN(n2123) );
  INV_X1 U1076 ( .A(n2123), .ZN(n756) );
  AOI21_X1 U1077 ( .B1(n2124), .B2(n757), .A(n756), .ZN(n758) );
  OAI21_X1 U1078 ( .B1(n760), .B2(n759), .A(n758), .ZN(n1872) );
  XNOR2_X1 U1079 ( .A(fmem_data[7]), .B(n1245), .ZN(n805) );
  OAI22_X1 U1080 ( .A1(n1251), .A2(n761), .B1(n1249), .B2(n805), .ZN(n794) );
  XNOR2_X1 U1081 ( .A(fmem_data[13]), .B(n849), .ZN(n790) );
  OAI22_X1 U1082 ( .A1(n875), .A2(n762), .B1(n871), .B2(n790), .ZN(n793) );
  NAND2_X1 U1083 ( .A1(n764), .A2(n763), .ZN(n1255) );
  BUF_X2 U1084 ( .A(n1255), .Z(n1512) );
  BUF_X4 U1085 ( .A(xmem_data[19]), .Z(n1324) );
  INV_X1 U1086 ( .A(n1324), .ZN(n766) );
  OR2_X1 U1087 ( .A1(n285), .A2(n766), .ZN(n765) );
  OAI22_X1 U1088 ( .A1(n1237), .A2(n766), .B1(n247), .B2(n765), .ZN(n792) );
  FA_X1 U1089 ( .A(n769), .B(n768), .CI(n767), .CO(n809), .S(n783) );
  XNOR2_X1 U1090 ( .A(n886), .B(fmem_data[9]), .ZN(n787) );
  OAI22_X1 U1091 ( .A1(n296), .A2(n770), .B1(n787), .B2(n1010), .ZN(n804) );
  XNOR2_X1 U1092 ( .A(n284), .B(n1324), .ZN(n771) );
  XNOR2_X1 U1093 ( .A(fmem_data[1]), .B(n1324), .ZN(n806) );
  OAI22_X1 U1094 ( .A1(n1237), .A2(n771), .B1(n247), .B2(n806), .ZN(n803) );
  XNOR2_X1 U1095 ( .A(fmem_data[5]), .B(n1269), .ZN(n807) );
  OAI22_X1 U1096 ( .A1(n723), .A2(n772), .B1(n1271), .B2(n807), .ZN(n802) );
  AOI21_X1 U1097 ( .B1(n774), .B2(n711), .A(n773), .ZN(n775) );
  INV_X1 U1098 ( .A(n775), .ZN(n786) );
  OR2_X1 U1099 ( .A1(n777), .A2(n776), .ZN(n785) );
  FA_X1 U1100 ( .A(n780), .B(n779), .CI(n778), .CO(n784), .S(n817) );
  FA_X1 U1101 ( .A(n783), .B(n782), .CI(n781), .CO(n827), .S(n837) );
  FA_X1 U1102 ( .A(n786), .B(n785), .CI(n784), .CO(n985), .S(n828) );
  XNOR2_X1 U1103 ( .A(n886), .B(fmem_data[10]), .ZN(n924) );
  OAI22_X1 U1104 ( .A1(n297), .A2(n787), .B1(n924), .B2(n1010), .ZN(n949) );
  BUF_X2 U1105 ( .A(n925), .Z(n1268) );
  XNOR2_X1 U1106 ( .A(n1266), .B(n229), .ZN(n797) );
  XNOR2_X1 U1107 ( .A(n1266), .B(fmem_data[4]), .ZN(n927) );
  BUF_X1 U1108 ( .A(n788), .Z(n1220) );
  OAI22_X1 U1109 ( .A1(n1268), .A2(n797), .B1(n927), .B2(n1220), .ZN(n948) );
  XNOR2_X1 U1110 ( .A(fmem_data[11]), .B(n890), .ZN(n795) );
  XNOR2_X1 U1111 ( .A(fmem_data[12]), .B(n890), .ZN(n930) );
  OAI22_X1 U1112 ( .A1(n1037), .A2(n795), .B1(n929), .B2(n930), .ZN(n947) );
  XNOR2_X1 U1113 ( .A(n4052), .B(n4064), .ZN(n900) );
  BUF_X2 U1114 ( .A(n900), .Z(n1584) );
  INV_X1 U1115 ( .A(n1584), .ZN(n789) );
  AND2_X1 U1116 ( .A1(n287), .A2(n789), .ZN(n860) );
  XNOR2_X1 U1117 ( .A(fmem_data[14]), .B(n849), .ZN(n874) );
  OAI22_X1 U1118 ( .A1(n875), .A2(n790), .B1(n871), .B2(n874), .ZN(n861) );
  XNOR2_X1 U1119 ( .A(n860), .B(n861), .ZN(n958) );
  XNOR2_X1 U1120 ( .A(fmem_data[31]), .B(n261), .ZN(n856) );
  XNOR2_X1 U1121 ( .A(n261), .B(fmem_data[15]), .ZN(n799) );
  OAI22_X1 U1122 ( .A1(n856), .A2(n857), .B1(n801), .B2(n799), .ZN(n957) );
  FA_X1 U1123 ( .A(n794), .B(n793), .CI(n792), .CO(n956), .S(n810) );
  OAI22_X1 U1124 ( .A1(n931), .A2(n796), .B1(n1036), .B2(n795), .ZN(n813) );
  OAI22_X1 U1125 ( .A1(n1356), .A2(n798), .B1(n797), .B2(n1353), .ZN(n812) );
  OAI22_X1 U1126 ( .A1(n801), .A2(n800), .B1(n799), .B2(n857), .ZN(n811) );
  FA_X1 U1127 ( .A(n804), .B(n803), .CI(n802), .CO(n954), .S(n808) );
  XNOR2_X1 U1128 ( .A(fmem_data[8]), .B(n1245), .ZN(n880) );
  OAI22_X1 U1129 ( .A1(n1251), .A2(n805), .B1(n1233), .B2(n880), .ZN(n864) );
  OAI22_X1 U1130 ( .A1(n1512), .A2(n806), .B1(n247), .B2(n878), .ZN(n863) );
  XNOR2_X1 U1131 ( .A(fmem_data[6]), .B(n1269), .ZN(n920) );
  OAI22_X1 U1132 ( .A1(n201), .A2(n807), .B1(n141), .B2(n920), .ZN(n862) );
  FA_X1 U1133 ( .A(n810), .B(n809), .CI(n808), .CO(n1055), .S(n829) );
  XNOR2_X1 U1134 ( .A(n1056), .B(n1055), .ZN(n820) );
  FA_X1 U1135 ( .A(n813), .B(n812), .CI(n811), .CO(n955), .S(n826) );
  FA_X1 U1136 ( .A(n816), .B(n815), .CI(n814), .CO(n825), .S(n822) );
  FA_X1 U1137 ( .A(n819), .B(n818), .CI(n817), .CO(n824), .S(n821) );
  FA_X1 U1138 ( .A(n823), .B(n822), .CI(n821), .CO(n832), .S(n833) );
  FA_X1 U1139 ( .A(n829), .B(n828), .CI(n827), .CO(n1070), .S(n830) );
  NOR2_X1 U1140 ( .A1(n1865), .A2(n1864), .ZN(n843) );
  FA_X1 U1141 ( .A(n832), .B(n831), .CI(n830), .CO(n1864), .S(n842) );
  NOR2_X1 U1142 ( .A1(n197), .A2(n841), .ZN(n1866) );
  NOR2_X1 U1143 ( .A1(n843), .A2(n1866), .ZN(n1852) );
  NAND2_X1 U1144 ( .A1(n842), .A2(n841), .ZN(n3676) );
  NAND2_X1 U1145 ( .A1(n1865), .A2(n1864), .ZN(n2148) );
  OAI21_X1 U1146 ( .B1(n843), .B2(n3676), .A(n2148), .ZN(n1855) );
  XNOR2_X1 U1147 ( .A(fmem_data[10]), .B(n252), .ZN(n851) );
  XNOR2_X1 U1148 ( .A(fmem_data[11]), .B(n252), .ZN(n888) );
  OAI22_X1 U1149 ( .A1(n1246), .A2(n851), .B1(n1249), .B2(n888), .ZN(n894) );
  XNOR2_X1 U1150 ( .A(fmem_data[4]), .B(n1324), .ZN(n854) );
  XNOR2_X1 U1151 ( .A(fmem_data[5]), .B(n1324), .ZN(n906) );
  OAI22_X1 U1152 ( .A1(n1237), .A2(n854), .B1(n247), .B2(n906), .ZN(n893) );
  XNOR2_X1 U1153 ( .A(n4062), .B(xmem_data[22]), .ZN(n844) );
  BUF_X4 U1154 ( .A(xmem_data[23]), .Z(n1610) );
  OR2_X1 U1155 ( .A1(n285), .A2(n213), .ZN(n845) );
  OAI22_X1 U1156 ( .A1(n1008), .A2(n213), .B1(n845), .B2(n1641), .ZN(n892) );
  XNOR2_X1 U1157 ( .A(n1231), .B(fmem_data[11]), .ZN(n923) );
  XNOR2_X1 U1158 ( .A(n1231), .B(fmem_data[12]), .ZN(n847) );
  OAI22_X1 U1159 ( .A1(n297), .A2(n923), .B1(n847), .B2(n1010), .ZN(n867) );
  XNOR2_X1 U1160 ( .A(xmem_data[21]), .B(n4052), .ZN(n846) );
  NAND2_X1 U1161 ( .A1(n900), .A2(n846), .ZN(n899) );
  BUF_X2 U1162 ( .A(n899), .Z(n1585) );
  BUF_X4 U1163 ( .A(xmem_data[21]), .Z(n1530) );
  XNOR2_X1 U1164 ( .A(fmem_data[1]), .B(n1530), .ZN(n921) );
  XNOR2_X1 U1165 ( .A(fmem_data[2]), .B(n1530), .ZN(n901) );
  OAI22_X1 U1166 ( .A1(n1585), .A2(n921), .B1(n1584), .B2(n901), .ZN(n866) );
  XNOR2_X1 U1167 ( .A(fmem_data[13]), .B(n890), .ZN(n928) );
  XNOR2_X1 U1168 ( .A(fmem_data[14]), .B(n189), .ZN(n848) );
  OAI22_X1 U1169 ( .A1(n1037), .A2(n928), .B1(n1036), .B2(n848), .ZN(n865) );
  XNOR2_X1 U1170 ( .A(n1231), .B(fmem_data[13]), .ZN(n887) );
  OAI22_X1 U1171 ( .A1(n296), .A2(n847), .B1(n887), .B2(n1010), .ZN(n904) );
  XNOR2_X1 U1172 ( .A(n1266), .B(fmem_data[6]), .ZN(n855) );
  XNOR2_X1 U1173 ( .A(n1266), .B(n238), .ZN(n905) );
  OAI22_X1 U1174 ( .A1(n1356), .A2(n855), .B1(n905), .B2(n1220), .ZN(n903) );
  XNOR2_X1 U1175 ( .A(fmem_data[15]), .B(n189), .ZN(n891) );
  OAI22_X1 U1176 ( .A1(n1037), .A2(n848), .B1(n929), .B2(n891), .ZN(n902) );
  XNOR2_X1 U1177 ( .A(fmem_data[31]), .B(n279), .ZN(n872) );
  AOI21_X1 U1178 ( .B1(n870), .B2(n871), .A(n872), .ZN(n850) );
  INV_X1 U1179 ( .A(n850), .ZN(n885) );
  XNOR2_X1 U1180 ( .A(fmem_data[9]), .B(n1245), .ZN(n879) );
  OAI22_X1 U1181 ( .A1(n1246), .A2(n879), .B1(n1233), .B2(n851), .ZN(n869) );
  INV_X1 U1182 ( .A(n1641), .ZN(n853) );
  AND2_X1 U1183 ( .A1(n285), .A2(n853), .ZN(n868) );
  OR2_X1 U1184 ( .A1(n869), .A2(n868), .ZN(n884) );
  XNOR2_X1 U1185 ( .A(fmem_data[7]), .B(n1269), .ZN(n919) );
  XNOR2_X1 U1186 ( .A(n258), .B(n1269), .ZN(n898) );
  OAI22_X1 U1187 ( .A1(n201), .A2(n919), .B1(n1271), .B2(n898), .ZN(n934) );
  OAI22_X1 U1188 ( .A1(n1237), .A2(n876), .B1(n1253), .B2(n854), .ZN(n933) );
  XNOR2_X1 U1189 ( .A(n1266), .B(fmem_data[5]), .ZN(n926) );
  OAI22_X1 U1190 ( .A1(n1268), .A2(n926), .B1(n855), .B2(n1353), .ZN(n932) );
  AOI21_X1 U1191 ( .B1(n858), .B2(n857), .A(n856), .ZN(n859) );
  INV_X1 U1192 ( .A(n859), .ZN(n979) );
  OR2_X1 U1193 ( .A1(n861), .A2(n860), .ZN(n978) );
  FA_X1 U1194 ( .A(n863), .B(n864), .CI(n862), .CO(n977), .S(n953) );
  FA_X1 U1195 ( .A(n867), .B(n866), .CI(n865), .CO(n910), .S(n989) );
  XNOR2_X1 U1196 ( .A(n869), .B(n868), .ZN(n914) );
  XNOR2_X1 U1197 ( .A(fmem_data[15]), .B(n849), .ZN(n873) );
  OAI22_X1 U1198 ( .A1(n872), .A2(n871), .B1(n870), .B2(n873), .ZN(n913) );
  OAI22_X1 U1199 ( .A1(n875), .A2(n874), .B1(n871), .B2(n873), .ZN(n946) );
  OR2_X1 U1200 ( .A1(n876), .A2(n249), .ZN(n877) );
  OAI21_X1 U1201 ( .B1(n1512), .B2(n878), .A(n877), .ZN(n945) );
  OAI22_X1 U1202 ( .A1(n1251), .A2(n880), .B1(n1249), .B2(n879), .ZN(n944) );
  OAI21_X1 U1203 ( .B1(n972), .B2(n971), .A(n973), .ZN(n882) );
  NAND2_X1 U1204 ( .A1(n972), .A2(n971), .ZN(n881) );
  NAND2_X1 U1205 ( .A1(n882), .A2(n881), .ZN(n1050) );
  FA_X1 U1206 ( .A(n885), .B(n884), .CI(n883), .CO(n1022), .S(n971) );
  XNOR2_X1 U1207 ( .A(n184), .B(n1269), .ZN(n897) );
  XNOR2_X1 U1208 ( .A(n203), .B(n1269), .ZN(n1012) );
  OAI22_X1 U1209 ( .A1(n723), .A2(n897), .B1(n1271), .B2(n1012), .ZN(n1030) );
  XNOR2_X1 U1210 ( .A(n1610), .B(fmem_data[1]), .ZN(n895) );
  XNOR2_X1 U1211 ( .A(n1610), .B(fmem_data[2]), .ZN(n1009) );
  OAI22_X1 U1212 ( .A1(n1008), .A2(n895), .B1(n1009), .B2(n1641), .ZN(n1029)
         );
  XNOR2_X1 U1213 ( .A(n886), .B(fmem_data[14]), .ZN(n1011) );
  OAI22_X1 U1214 ( .A1(n297), .A2(n887), .B1(n1011), .B2(n1010), .ZN(n1028) );
  XNOR2_X1 U1215 ( .A(fmem_data[12]), .B(n252), .ZN(n1023) );
  OAI22_X1 U1216 ( .A1(n1246), .A2(n888), .B1(n1233), .B2(n1023), .ZN(n1040)
         );
  INV_X1 U1217 ( .A(n191), .ZN(n889) );
  AND2_X1 U1218 ( .A1(n285), .A2(n889), .ZN(n1039) );
  XNOR2_X1 U1219 ( .A(n1040), .B(n1039), .ZN(n1007) );
  XNOR2_X1 U1220 ( .A(fmem_data[31]), .B(n189), .ZN(n1035) );
  OAI22_X1 U1221 ( .A1(n1035), .A2(n929), .B1(n1037), .B2(n891), .ZN(n1006) );
  FA_X1 U1222 ( .A(n894), .B(n893), .CI(n892), .CO(n1005), .S(n911) );
  XNOR2_X1 U1223 ( .A(n1050), .B(n1049), .ZN(n939) );
  XNOR2_X1 U1224 ( .A(n1610), .B(n286), .ZN(n896) );
  OAI22_X1 U1225 ( .A1(n1008), .A2(n896), .B1(n895), .B2(n1641), .ZN(n917) );
  OAI22_X1 U1226 ( .A1(n723), .A2(n898), .B1(n219), .B2(n897), .ZN(n916) );
  XNOR2_X1 U1227 ( .A(n229), .B(n1530), .ZN(n907) );
  OAI22_X1 U1228 ( .A1(n1585), .A2(n901), .B1(n1533), .B2(n907), .ZN(n915) );
  FA_X1 U1229 ( .A(n904), .B(n903), .CI(n902), .CO(n1015), .S(n909) );
  XNOR2_X1 U1230 ( .A(n1016), .B(n1015), .ZN(n908) );
  XNOR2_X1 U1231 ( .A(n1266), .B(fmem_data[8]), .ZN(n1031) );
  OAI22_X1 U1232 ( .A1(n1356), .A2(n905), .B1(n1031), .B2(n1353), .ZN(n1043)
         );
  XNOR2_X1 U1233 ( .A(n4063), .B(n300), .ZN(n1024) );
  OAI22_X1 U1234 ( .A1(n1237), .A2(n906), .B1(n1253), .B2(n1024), .ZN(n1042)
         );
  XNOR2_X1 U1235 ( .A(fmem_data[4]), .B(n1530), .ZN(n1034) );
  OAI22_X1 U1236 ( .A1(n1585), .A2(n907), .B1(n1584), .B2(n1034), .ZN(n1041)
         );
  XNOR2_X1 U1237 ( .A(n908), .B(n1014), .ZN(n1001) );
  FA_X1 U1238 ( .A(n911), .B(n910), .CI(n909), .CO(n1000), .S(n972) );
  XNOR2_X1 U1239 ( .A(n1001), .B(n1000), .ZN(n938) );
  FA_X1 U1240 ( .A(n914), .B(n913), .CI(n912), .CO(n970), .S(n988) );
  FA_X1 U1241 ( .A(n917), .B(n916), .CI(n915), .CO(n1016), .S(n969) );
  OR2_X1 U1242 ( .A1(n287), .A2(n206), .ZN(n918) );
  OAI22_X1 U1243 ( .A1(n1532), .A2(n206), .B1(n1533), .B2(n918), .ZN(n961) );
  OAI22_X1 U1244 ( .A1(n201), .A2(n920), .B1(n1271), .B2(n919), .ZN(n960) );
  XNOR2_X1 U1245 ( .A(n287), .B(n1530), .ZN(n922) );
  OAI22_X1 U1246 ( .A1(n1585), .A2(n922), .B1(n1533), .B2(n921), .ZN(n959) );
  OAI22_X1 U1247 ( .A1(n295), .A2(n924), .B1(n923), .B2(n1010), .ZN(n952) );
  OAI22_X1 U1248 ( .A1(n1356), .A2(n927), .B1(n926), .B2(n1220), .ZN(n951) );
  OAI22_X1 U1249 ( .A1(n931), .A2(n930), .B1(n929), .B2(n928), .ZN(n950) );
  NAND2_X1 U1250 ( .A1(n940), .A2(n941), .ZN(n937) );
  FA_X1 U1251 ( .A(n934), .B(n933), .CI(n932), .CO(n883), .S(n942) );
  OR2_X1 U1252 ( .A1(n940), .A2(n941), .ZN(n935) );
  NAND2_X1 U1253 ( .A1(n942), .A2(n935), .ZN(n936) );
  NAND2_X1 U1254 ( .A1(n937), .A2(n936), .ZN(n968) );
  XNOR2_X1 U1255 ( .A(n941), .B(n940), .ZN(n943) );
  XNOR2_X1 U1256 ( .A(n943), .B(n942), .ZN(n992) );
  FA_X1 U1257 ( .A(n946), .B(n945), .CI(n944), .CO(n912), .S(n982) );
  FA_X1 U1258 ( .A(n949), .B(n948), .CI(n947), .CO(n981), .S(n984) );
  FA_X1 U1259 ( .A(n952), .B(n951), .CI(n950), .CO(n941), .S(n980) );
  OR2_X1 U1260 ( .A1(n992), .A2(n991), .ZN(n965) );
  FA_X1 U1261 ( .A(n955), .B(n954), .CI(n953), .CO(n1064), .S(n1056) );
  FA_X1 U1262 ( .A(n958), .B(n957), .CI(n956), .CO(n1062), .S(n983) );
  FA_X1 U1263 ( .A(n961), .B(n960), .CI(n959), .CO(n940), .S(n1061) );
  NAND2_X1 U1264 ( .A1(n1064), .A2(n962), .ZN(n964) );
  NAND2_X1 U1265 ( .A1(n964), .A2(n963), .ZN(n993) );
  NAND2_X1 U1266 ( .A1(n992), .A2(n991), .ZN(n966) );
  FA_X1 U1267 ( .A(n970), .B(n969), .CI(n968), .CO(n999), .S(n995) );
  NOR2_X2 U1268 ( .A1(n1085), .A2(n1084), .ZN(n1879) );
  FA_X1 U1269 ( .A(n979), .B(n978), .CI(n977), .CO(n990), .S(n1065) );
  FA_X1 U1270 ( .A(n982), .B(n981), .CI(n980), .CO(n991), .S(n1066) );
  FA_X1 U1271 ( .A(n985), .B(n984), .CI(n983), .CO(n1067), .S(n1069) );
  FA_X1 U1272 ( .A(n990), .B(n989), .CI(n988), .CO(n973), .S(n1072) );
  XNOR2_X1 U1273 ( .A(n992), .B(n991), .ZN(n994) );
  XNOR2_X1 U1274 ( .A(n994), .B(n993), .ZN(n1071) );
  XNOR2_X1 U1275 ( .A(n996), .B(n995), .ZN(n998) );
  XNOR2_X1 U1276 ( .A(n998), .B(n997), .ZN(n1083) );
  NOR2_X1 U1277 ( .A1(n1082), .A2(n1083), .ZN(n3660) );
  NOR2_X1 U1278 ( .A1(n1879), .A2(n3660), .ZN(n2028) );
  INV_X1 U1279 ( .A(n999), .ZN(n1004) );
  FA_X1 U1280 ( .A(n1007), .B(n1006), .CI(n1005), .CO(n1387), .S(n1020) );
  XNOR2_X1 U1281 ( .A(n1610), .B(n228), .ZN(n1358) );
  OAI22_X1 U1282 ( .A1(n1008), .A2(n1009), .B1(n1358), .B2(n1641), .ZN(n1388)
         );
  XNOR2_X1 U1283 ( .A(n1231), .B(fmem_data[15]), .ZN(n1370) );
  OAI22_X1 U1284 ( .A1(n297), .A2(n1011), .B1(n1370), .B2(n1010), .ZN(n1390)
         );
  XNOR2_X1 U1285 ( .A(fmem_data[11]), .B(n1113), .ZN(n1360) );
  OAI22_X1 U1286 ( .A1(n201), .A2(n1012), .B1(n219), .B2(n1360), .ZN(n1389) );
  XOR2_X1 U1287 ( .A(n1390), .B(n1389), .Z(n1013) );
  XOR2_X1 U1288 ( .A(n1388), .B(n1013), .Z(n1386) );
  FA_X1 U1289 ( .A(n1022), .B(n1021), .CI(n1020), .CO(n1424), .S(n1049) );
  XNOR2_X1 U1290 ( .A(fmem_data[13]), .B(n252), .ZN(n1234) );
  OAI22_X1 U1291 ( .A1(n1251), .A2(n1023), .B1(n1234), .B2(n1233), .ZN(n1375)
         );
  OAI22_X1 U1292 ( .A1(n1512), .A2(n1024), .B1(n1236), .B2(n247), .ZN(n1374)
         );
  XNOR2_X1 U1293 ( .A(xmem_data[25]), .B(n313), .ZN(n1025) );
  INV_X1 U1294 ( .A(n244), .ZN(n1027) );
  OR2_X1 U1295 ( .A1(n287), .A2(n1027), .ZN(n1026) );
  OAI22_X1 U1296 ( .A1(n274), .A2(n1027), .B1(n191), .B2(n1026), .ZN(n1373) );
  FA_X1 U1297 ( .A(n1030), .B(n1029), .CI(n1028), .CO(n1402), .S(n1021) );
  XNOR2_X1 U1298 ( .A(n1266), .B(fmem_data[9]), .ZN(n1355) );
  OAI22_X1 U1299 ( .A1(n1268), .A2(n1031), .B1(n1355), .B2(n1220), .ZN(n1396)
         );
  XNOR2_X1 U1300 ( .A(n285), .B(n245), .ZN(n1033) );
  OAI22_X1 U1301 ( .A1(n196), .A2(n1033), .B1(n140), .B2(n1238), .ZN(n1395) );
  XNOR2_X1 U1302 ( .A(fmem_data[5]), .B(n1530), .ZN(n1239) );
  OAI22_X1 U1303 ( .A1(n1532), .A2(n1034), .B1(n1584), .B2(n1239), .ZN(n1394)
         );
  AOI21_X1 U1304 ( .B1(n1037), .B2(n1036), .A(n1035), .ZN(n1038) );
  INV_X1 U1305 ( .A(n1038), .ZN(n1378) );
  OR2_X1 U1306 ( .A1(n1040), .A2(n1039), .ZN(n1377) );
  FA_X1 U1307 ( .A(n1043), .B(n1042), .CI(n1041), .CO(n1376), .S(n1014) );
  XNOR2_X1 U1308 ( .A(n1427), .B(n1426), .ZN(n1044) );
  XNOR2_X1 U1309 ( .A(n1424), .B(n1044), .ZN(n1463) );
  INV_X1 U1310 ( .A(n1050), .ZN(n1046) );
  NAND2_X1 U1311 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  OR2_X2 U1312 ( .A1(n1087), .A2(n1086), .ZN(n1874) );
  INV_X1 U1313 ( .A(n1056), .ZN(n1054) );
  INV_X1 U1314 ( .A(n1055), .ZN(n1053) );
  NAND2_X1 U1315 ( .A1(n1054), .A2(n1053), .ZN(n1058) );
  AND2_X1 U1316 ( .A1(n1056), .A2(n1055), .ZN(n1057) );
  AOI21_X1 U1317 ( .B1(n1059), .B2(n1058), .A(n1057), .ZN(n1060) );
  INV_X1 U1318 ( .A(n1060), .ZN(n1076) );
  XNOR2_X1 U1319 ( .A(n1066), .B(n1065), .ZN(n1068) );
  XNOR2_X1 U1320 ( .A(n1068), .B(n1067), .ZN(n1074) );
  FA_X1 U1321 ( .A(n1073), .B(n1072), .CI(n1071), .CO(n1082), .S(n1081) );
  FA_X1 U1322 ( .A(n1076), .B(n1075), .CI(n1074), .CO(n1080), .S(n1079) );
  NAND2_X1 U1323 ( .A1(n2075), .A2(n2133), .ZN(n1869) );
  INV_X1 U1324 ( .A(n208), .ZN(n1077) );
  NAND2_X1 U1325 ( .A1(n336), .A2(n1077), .ZN(n1092) );
  AOI21_X1 U1326 ( .B1(n2076), .B2(n2133), .A(n217), .ZN(n1868) );
  NAND2_X1 U1327 ( .A1(n1083), .A2(n1082), .ZN(n3670) );
  OAI21_X1 U1328 ( .B1(n1868), .B2(n3660), .A(n3670), .ZN(n1090) );
  NOR2_X1 U1329 ( .A1(n1879), .A2(n2027), .ZN(n1089) );
  NAND2_X1 U1330 ( .A1(n1085), .A2(n1084), .ZN(n3663) );
  NAND2_X1 U1331 ( .A1(n1087), .A2(n1086), .ZN(n2029) );
  OAI21_X1 U1332 ( .B1(n210), .B2(n3663), .A(n185), .ZN(n1088) );
  AOI21_X1 U1333 ( .B1(n1090), .B2(n1089), .A(n1088), .ZN(n1091) );
  OAI21_X1 U1334 ( .B1(n2131), .B2(n1092), .A(n1091), .ZN(n2175) );
  INV_X1 U1335 ( .A(n2175), .ZN(n1826) );
  XNOR2_X1 U1336 ( .A(n1610), .B(n258), .ZN(n1118) );
  XNOR2_X1 U1337 ( .A(n1610), .B(fmem_data[9]), .ZN(n1154) );
  OAI22_X1 U1338 ( .A1(n1008), .A2(n1118), .B1(n1154), .B2(n1641), .ZN(n1109)
         );
  XNOR2_X1 U1339 ( .A(n4054), .B(xmem_data[30]), .ZN(n1093) );
  XNOR2_X1 U1340 ( .A(xmem_data[29]), .B(xmem_data[30]), .ZN(n1123) );
  NAND2_X1 U1341 ( .A1(n1093), .A2(n1123), .ZN(n1571) );
  XNOR2_X1 U1342 ( .A(xmem_data[31]), .B(n287), .ZN(n1094) );
  XNOR2_X1 U1343 ( .A(xmem_data[31]), .B(fmem_data[1]), .ZN(n1099) );
  OAI22_X1 U1344 ( .A1(n1547), .A2(n1094), .B1(n1099), .B2(n1743), .ZN(n1108)
         );
  XOR2_X1 U1345 ( .A(n4065), .B(n4066), .Z(n1235) );
  NAND2_X1 U1346 ( .A1(n1095), .A2(n1696), .ZN(n1104) );
  BUF_X2 U1347 ( .A(n1104), .Z(n1312) );
  BUF_X4 U1348 ( .A(n1096), .Z(n1693) );
  XNOR2_X1 U1349 ( .A(fmem_data[4]), .B(n1693), .ZN(n1105) );
  OR2_X1 U1350 ( .A1(n1159), .A2(n307), .ZN(n1097) );
  OAI21_X1 U1351 ( .B1(n1312), .B2(n1105), .A(n1097), .ZN(n1107) );
  XNOR2_X1 U1352 ( .A(fmem_data[10]), .B(n1530), .ZN(n1103) );
  XNOR2_X1 U1353 ( .A(fmem_data[11]), .B(n1530), .ZN(n1145) );
  OAI22_X1 U1354 ( .A1(n1532), .A2(n1103), .B1(n1533), .B2(n1145), .ZN(n1134)
         );
  OR2_X1 U1355 ( .A1(n285), .A2(n4054), .ZN(n1098) );
  OAI22_X1 U1356 ( .A1(n1747), .A2(n4054), .B1(n1098), .B2(n1743), .ZN(n1133)
         );
  XNOR2_X1 U1357 ( .A(n1266), .B(fmem_data[14]), .ZN(n1106) );
  XNOR2_X1 U1358 ( .A(n1266), .B(fmem_data[15]), .ZN(n1144) );
  OAI22_X1 U1359 ( .A1(n1356), .A2(n1106), .B1(n1144), .B2(n1220), .ZN(n1132)
         );
  XNOR2_X1 U1360 ( .A(fmem_data[13]), .B(n1324), .ZN(n1102) );
  XNOR2_X1 U1361 ( .A(fmem_data[14]), .B(n1324), .ZN(n1164) );
  OAI22_X1 U1362 ( .A1(n1237), .A2(n1102), .B1(n1253), .B2(n1164), .ZN(n1162)
         );
  XNOR2_X1 U1363 ( .A(fmem_data[7]), .B(n246), .ZN(n1100) );
  XNOR2_X1 U1364 ( .A(n182), .B(fmem_data[8]), .ZN(n1163) );
  OAI22_X1 U1365 ( .A1(n196), .A2(n1100), .B1(n191), .B2(n1163), .ZN(n1161) );
  XNOR2_X1 U1366 ( .A(xmem_data[31]), .B(fmem_data[2]), .ZN(n1139) );
  OAI22_X1 U1367 ( .A1(n1571), .A2(n1099), .B1(n1139), .B2(n1743), .ZN(n1160)
         );
  XNOR2_X1 U1368 ( .A(n245), .B(fmem_data[6]), .ZN(n1116) );
  OAI22_X1 U1369 ( .A1(n274), .A2(n1116), .B1(n191), .B2(n1100), .ZN(n1143) );
  XNOR2_X1 U1370 ( .A(xmem_data[27]), .B(xmem_data[28]), .ZN(n1128) );
  NAND2_X1 U1371 ( .A1(n1128), .A2(n1101), .ZN(n1127) );
  XNOR2_X1 U1372 ( .A(fmem_data[2]), .B(n1711), .ZN(n1122) );
  BUF_X2 U1373 ( .A(n1128), .Z(n1731) );
  OAI22_X1 U1374 ( .A1(n1713), .A2(n1122), .B1(n1156), .B2(n1731), .ZN(n1142)
         );
  XNOR2_X1 U1375 ( .A(n4056), .B(n300), .ZN(n1117) );
  OAI22_X1 U1376 ( .A1(n1237), .A2(n1117), .B1(n247), .B2(n1102), .ZN(n1141)
         );
  XNOR2_X1 U1377 ( .A(fmem_data[9]), .B(n1530), .ZN(n1114) );
  OAI22_X1 U1378 ( .A1(n1585), .A2(n1114), .B1(n1533), .B2(n1103), .ZN(n1203)
         );
  BUF_X2 U1379 ( .A(n1104), .Z(n1697) );
  XNOR2_X1 U1380 ( .A(n1638), .B(n229), .ZN(n1111) );
  OAI22_X1 U1381 ( .A1(n1697), .A2(n1111), .B1(n306), .B2(n1105), .ZN(n1202)
         );
  XNOR2_X1 U1382 ( .A(n1266), .B(fmem_data[13]), .ZN(n1110) );
  OAI22_X1 U1383 ( .A1(n1268), .A2(n1110), .B1(n1106), .B2(n1353), .ZN(n1201)
         );
  FA_X1 U1384 ( .A(n1108), .B(n1109), .CI(n1107), .CO(n1167), .S(n1185) );
  XNOR2_X1 U1385 ( .A(n1266), .B(fmem_data[12]), .ZN(n1221) );
  OAI22_X1 U1386 ( .A1(n1356), .A2(n1221), .B1(n1110), .B2(n1220), .ZN(n1263)
         );
  XNOR2_X1 U1387 ( .A(fmem_data[2]), .B(n1693), .ZN(n1222) );
  OR2_X1 U1388 ( .A1(n1111), .A2(n306), .ZN(n1112) );
  OAI21_X1 U1389 ( .B1(n1312), .B2(n1222), .A(n1112), .ZN(n1262) );
  XNOR2_X1 U1390 ( .A(fmem_data[14]), .B(n1113), .ZN(n1223) );
  XNOR2_X1 U1391 ( .A(fmem_data[15]), .B(n1269), .ZN(n1125) );
  OAI22_X1 U1392 ( .A1(n723), .A2(n1223), .B1(n141), .B2(n1125), .ZN(n1261) );
  OAI22_X1 U1393 ( .A1(n1585), .A2(n1197), .B1(n1584), .B2(n1114), .ZN(n1227)
         );
  OR2_X1 U1394 ( .A1(n286), .A2(n331), .ZN(n1115) );
  OAI22_X1 U1395 ( .A1(n1713), .A2(n331), .B1(n1115), .B2(n1731), .ZN(n1226)
         );
  XNOR2_X1 U1396 ( .A(n1610), .B(fmem_data[6]), .ZN(n1194) );
  XNOR2_X1 U1397 ( .A(n1610), .B(fmem_data[7]), .ZN(n1120) );
  OAI22_X1 U1398 ( .A1(n1008), .A2(n1194), .B1(n1120), .B2(n1641), .ZN(n1225)
         );
  XNOR2_X1 U1399 ( .A(n182), .B(fmem_data[5]), .ZN(n1126) );
  OAI22_X1 U1400 ( .A1(n276), .A2(n1126), .B1(n191), .B2(n1116), .ZN(n1174) );
  XNOR2_X1 U1401 ( .A(fmem_data[11]), .B(n1324), .ZN(n1131) );
  OAI22_X1 U1402 ( .A1(n1237), .A2(n1131), .B1(n1253), .B2(n1117), .ZN(n1173)
         );
  XNOR2_X1 U1403 ( .A(n1174), .B(n1173), .ZN(n1121) );
  OR2_X1 U1404 ( .A1(n1118), .A2(n1641), .ZN(n1119) );
  XNOR2_X1 U1405 ( .A(n1121), .B(n1172), .ZN(n1283) );
  XNOR2_X1 U1406 ( .A(fmem_data[1]), .B(n281), .ZN(n1129) );
  OAI22_X1 U1407 ( .A1(n1713), .A2(n1129), .B1(n1122), .B2(n1731), .ZN(n1171)
         );
  INV_X1 U1408 ( .A(n231), .ZN(n1124) );
  AND2_X1 U1409 ( .A1(n285), .A2(n1124), .ZN(n1170) );
  XNOR2_X1 U1410 ( .A(n1171), .B(n1170), .ZN(n1206) );
  XNOR2_X1 U1411 ( .A(fmem_data[31]), .B(n1113), .ZN(n1168) );
  OAI22_X1 U1412 ( .A1(n1168), .A2(n219), .B1(n201), .B2(n1125), .ZN(n1205) );
  XNOR2_X1 U1413 ( .A(fmem_data[4]), .B(n246), .ZN(n1196) );
  OAI22_X1 U1414 ( .A1(n276), .A2(n1196), .B1(n140), .B2(n1126), .ZN(n1219) );
  XNOR2_X1 U1415 ( .A(n284), .B(n281), .ZN(n1130) );
  OAI22_X1 U1416 ( .A1(n1732), .A2(n1130), .B1(n1129), .B2(n1731), .ZN(n1218)
         );
  OAI22_X1 U1417 ( .A1(n1512), .A2(n1192), .B1(n247), .B2(n1131), .ZN(n1217)
         );
  FA_X1 U1418 ( .A(n1134), .B(n1132), .CI(n1133), .CO(n1166), .S(n1298) );
  INV_X1 U1419 ( .A(n1298), .ZN(n1135) );
  XNOR2_X1 U1420 ( .A(xmem_data[31]), .B(n228), .ZN(n1308) );
  OAI22_X1 U1421 ( .A1(n1547), .A2(n1139), .B1(n1308), .B2(n1743), .ZN(n1328)
         );
  XNOR2_X1 U1422 ( .A(fmem_data[4]), .B(n281), .ZN(n1155) );
  XNOR2_X1 U1423 ( .A(fmem_data[5]), .B(n281), .ZN(n1316) );
  OAI22_X1 U1424 ( .A1(n1713), .A2(n1155), .B1(n1316), .B2(n1731), .ZN(n1327)
         );
  XNOR2_X1 U1425 ( .A(fmem_data[6]), .B(n1638), .ZN(n1157) );
  OR2_X1 U1426 ( .A1(n1311), .A2(n307), .ZN(n1140) );
  OAI21_X1 U1427 ( .B1(n1312), .B2(n1157), .A(n1140), .ZN(n1326) );
  FA_X1 U1428 ( .A(n1141), .B(n1143), .CI(n1142), .CO(n1180), .S(n1187) );
  XNOR2_X1 U1429 ( .A(fmem_data[31]), .B(n1266), .ZN(n1150) );
  OAI22_X1 U1430 ( .A1(n1150), .A2(n1353), .B1(n1268), .B2(n1144), .ZN(n1178)
         );
  XNOR2_X1 U1431 ( .A(fmem_data[12]), .B(n1530), .ZN(n1149) );
  OAI22_X1 U1432 ( .A1(n1585), .A2(n1145), .B1(n1584), .B2(n1149), .ZN(n1177)
         );
  NAND2_X1 U1433 ( .A1(n1180), .A2(n1146), .ZN(n1148) );
  NAND2_X1 U1434 ( .A1(n1148), .A2(n1147), .ZN(n1333) );
  XNOR2_X1 U1435 ( .A(fmem_data[13]), .B(n1530), .ZN(n1317) );
  OAI22_X1 U1436 ( .A1(n1585), .A2(n1149), .B1(n1533), .B2(n1317), .ZN(n1315)
         );
  XNOR2_X1 U1437 ( .A(n1610), .B(n203), .ZN(n1153) );
  XNOR2_X1 U1438 ( .A(n1610), .B(fmem_data[11]), .ZN(n1319) );
  OAI22_X1 U1439 ( .A1(n1008), .A2(n1153), .B1(n1319), .B2(n1641), .ZN(n1314)
         );
  AOI21_X1 U1440 ( .B1(n1268), .B2(n1353), .A(n1150), .ZN(n1151) );
  INV_X1 U1441 ( .A(n1151), .ZN(n1313) );
  XNOR2_X1 U1442 ( .A(n1152), .B(n1332), .ZN(n1338) );
  XNOR2_X1 U1443 ( .A(n1339), .B(n1338), .ZN(n1184) );
  OAI22_X1 U1444 ( .A1(n1008), .A2(n1154), .B1(n1153), .B2(n1641), .ZN(n1183)
         );
  OAI22_X1 U1445 ( .A1(n1732), .A2(n1156), .B1(n1155), .B2(n1731), .ZN(n1322)
         );
  INV_X1 U1446 ( .A(n1322), .ZN(n1182) );
  OR2_X1 U1447 ( .A1(n1157), .A2(n307), .ZN(n1158) );
  OAI21_X1 U1448 ( .B1(n1312), .B2(n1159), .A(n1158), .ZN(n1181) );
  FA_X1 U1449 ( .A(n1162), .B(n1161), .CI(n1160), .CO(n1330), .S(n1165) );
  XNOR2_X1 U1450 ( .A(n182), .B(fmem_data[9]), .ZN(n1309) );
  OAI22_X1 U1451 ( .A1(n276), .A2(n1163), .B1(n140), .B2(n1309), .ZN(n1323) );
  XNOR2_X1 U1452 ( .A(fmem_data[15]), .B(n1324), .ZN(n1325) );
  OAI22_X1 U1453 ( .A1(n1237), .A2(n1164), .B1(n1253), .B2(n1325), .ZN(n1321)
         );
  FA_X1 U1454 ( .A(n1167), .B(n1166), .CI(n1165), .CO(n1306), .S(n1210) );
  AOI21_X1 U1455 ( .B1(n201), .B2(n1271), .A(n1168), .ZN(n1169) );
  INV_X1 U1456 ( .A(n1169), .ZN(n1190) );
  OR2_X1 U1457 ( .A1(n1171), .A2(n1170), .ZN(n1189) );
  OAI21_X1 U1458 ( .B1(n1173), .B2(n1174), .A(n1172), .ZN(n1176) );
  NAND2_X1 U1459 ( .A1(n1174), .A2(n1173), .ZN(n1175) );
  NAND2_X1 U1460 ( .A1(n1176), .A2(n1175), .ZN(n1188) );
  XNOR2_X1 U1461 ( .A(n1178), .B(n1177), .ZN(n1179) );
  XNOR2_X1 U1462 ( .A(n1180), .B(n1179), .ZN(n1208) );
  FA_X1 U1463 ( .A(n1183), .B(n1182), .CI(n1181), .CO(n1331), .S(n1207) );
  FA_X1 U1464 ( .A(n1187), .B(n1186), .CI(n1185), .CO(n1211), .S(n1304) );
  FA_X1 U1465 ( .A(n1190), .B(n1189), .CI(n1188), .CO(n1209), .S(n1303) );
  XNOR2_X1 U1466 ( .A(fmem_data[31]), .B(n252), .ZN(n1247) );
  AOI21_X1 U1467 ( .B1(n1246), .B2(n1233), .A(n1247), .ZN(n1191) );
  INV_X1 U1468 ( .A(n1191), .ZN(n1230) );
  XNOR2_X1 U1469 ( .A(n4057), .B(n300), .ZN(n1252) );
  OAI22_X1 U1470 ( .A1(n1512), .A2(n1252), .B1(n1253), .B2(n1192), .ZN(n1244)
         );
  INV_X1 U1471 ( .A(n1731), .ZN(n1193) );
  AND2_X1 U1472 ( .A1(n1193), .A2(n286), .ZN(n1243) );
  OR2_X1 U1473 ( .A1(n1244), .A2(n1243), .ZN(n1229) );
  XNOR2_X1 U1474 ( .A(n1610), .B(fmem_data[5]), .ZN(n1264) );
  OR2_X1 U1475 ( .A1(n1194), .A2(n1641), .ZN(n1195) );
  OAI21_X1 U1476 ( .B1(n1008), .B2(n1264), .A(n1195), .ZN(n1281) );
  XNOR2_X1 U1477 ( .A(n245), .B(n227), .ZN(n1256) );
  OAI22_X1 U1478 ( .A1(n275), .A2(n1256), .B1(n140), .B2(n1196), .ZN(n1280) );
  OAI22_X1 U1479 ( .A1(n1532), .A2(n1275), .B1(n1584), .B2(n1197), .ZN(n1279)
         );
  OR2_X1 U1480 ( .A1(n1279), .A2(n1280), .ZN(n1198) );
  NAND2_X1 U1481 ( .A1(n1281), .A2(n1198), .ZN(n1200) );
  NAND2_X1 U1482 ( .A1(n1280), .A2(n1279), .ZN(n1199) );
  NAND2_X1 U1483 ( .A1(n1200), .A2(n1199), .ZN(n1228) );
  FA_X1 U1484 ( .A(n1203), .B(n1202), .CI(n1201), .CO(n1186), .S(n1215) );
  FA_X1 U1485 ( .A(n1206), .B(n1205), .CI(n1204), .CO(n1299), .S(n1214) );
  FA_X1 U1486 ( .A(n1208), .B(n1207), .CI(n1209), .CO(n1305), .S(n1344) );
  XNOR2_X1 U1487 ( .A(n1210), .B(n1211), .ZN(n1212) );
  XNOR2_X1 U1488 ( .A(n1213), .B(n1212), .ZN(n1343) );
  XNOR2_X1 U1489 ( .A(n288), .B(n1900), .ZN(n1809) );
  FA_X1 U1490 ( .A(n1216), .B(n1215), .CI(n1214), .CO(n1302), .S(n1467) );
  FA_X1 U1491 ( .A(n1219), .B(n1217), .CI(n1218), .CO(n1204), .S(n1288) );
  XNOR2_X1 U1492 ( .A(n1266), .B(fmem_data[11]), .ZN(n1267) );
  OAI22_X1 U1493 ( .A1(n1268), .A2(n1267), .B1(n1221), .B2(n1220), .ZN(n1242)
         );
  XNOR2_X1 U1494 ( .A(fmem_data[1]), .B(n1693), .ZN(n1277) );
  OAI22_X1 U1495 ( .A1(n1312), .A2(n1277), .B1(n306), .B2(n1222), .ZN(n1241)
         );
  XNOR2_X1 U1496 ( .A(fmem_data[13]), .B(n1269), .ZN(n1270) );
  OAI22_X1 U1497 ( .A1(n201), .A2(n1270), .B1(n1271), .B2(n1223), .ZN(n1240)
         );
  FA_X1 U1498 ( .A(n1227), .B(n1226), .CI(n1225), .CO(n1284), .S(n1286) );
  FA_X1 U1499 ( .A(n1230), .B(n1229), .CI(n1228), .CO(n1216), .S(n1478) );
  XNOR2_X1 U1500 ( .A(fmem_data[31]), .B(n1231), .ZN(n1372) );
  AOI21_X1 U1501 ( .B1(n1010), .B2(n296), .A(n1372), .ZN(n1232) );
  INV_X1 U1502 ( .A(n1232), .ZN(n1367) );
  OAI22_X1 U1503 ( .A1(n1246), .A2(n1234), .B1(n1233), .B2(n1250), .ZN(n1369)
         );
  AND2_X1 U1504 ( .A1(n287), .A2(n305), .ZN(n1368) );
  OR2_X1 U1505 ( .A1(n1369), .A2(n1368), .ZN(n1366) );
  XOR2_X1 U1506 ( .A(fmem_data[8]), .B(n300), .Z(n1254) );
  OAI22_X1 U1507 ( .A1(n1512), .A2(n1236), .B1(n1253), .B2(n1254), .ZN(n1399)
         );
  OAI22_X1 U1508 ( .A1(n275), .A2(n1238), .B1(n140), .B2(n1257), .ZN(n1398) );
  XNOR2_X1 U1509 ( .A(fmem_data[6]), .B(n1530), .ZN(n1276) );
  OAI22_X1 U1510 ( .A1(n1532), .A2(n1239), .B1(n1584), .B2(n1276), .ZN(n1397)
         );
  FA_X1 U1511 ( .A(n1242), .B(n1240), .CI(n1241), .CO(n1287), .S(n1441) );
  XNOR2_X1 U1512 ( .A(n1243), .B(n1244), .ZN(n1260) );
  OAI22_X1 U1513 ( .A1(n1247), .A2(n1249), .B1(n1246), .B2(n1248), .ZN(n1259)
         );
  OAI22_X1 U1514 ( .A1(n1251), .A2(n1250), .B1(n1249), .B2(n1248), .ZN(n1352)
         );
  OAI22_X1 U1515 ( .A1(n1237), .A2(n1254), .B1(n1253), .B2(n1252), .ZN(n1351)
         );
  OAI22_X1 U1516 ( .A1(n1257), .A2(n275), .B1(n140), .B2(n1256), .ZN(n1350) );
  FA_X1 U1517 ( .A(n1259), .B(n1260), .CI(n1258), .CO(n1476), .S(n1440) );
  XNOR2_X1 U1518 ( .A(n1610), .B(n233), .ZN(n1357) );
  OR2_X1 U1519 ( .A1(n1264), .A2(n1641), .ZN(n1265) );
  OAI21_X1 U1520 ( .B1(n1008), .B2(n1357), .A(n1265), .ZN(n1363) );
  XNOR2_X1 U1521 ( .A(n1266), .B(fmem_data[10]), .ZN(n1354) );
  OAI22_X1 U1522 ( .A1(n1268), .A2(n1354), .B1(n1267), .B2(n1353), .ZN(n1361)
         );
  XNOR2_X1 U1523 ( .A(fmem_data[12]), .B(n1269), .ZN(n1359) );
  OAI22_X1 U1524 ( .A1(n723), .A2(n1359), .B1(n141), .B2(n1270), .ZN(n1362) );
  OAI21_X1 U1525 ( .B1(n1363), .B2(n1361), .A(n1362), .ZN(n1273) );
  NAND2_X1 U1526 ( .A1(n1363), .A2(n1361), .ZN(n1272) );
  NAND2_X1 U1527 ( .A1(n1273), .A2(n1272), .ZN(n1445) );
  OR2_X1 U1528 ( .A1(n284), .A2(n312), .ZN(n1274) );
  OAI22_X1 U1529 ( .A1(n1312), .A2(n312), .B1(n307), .B2(n1274), .ZN(n1412) );
  OAI22_X1 U1530 ( .A1(n1585), .A2(n1276), .B1(n1584), .B2(n1275), .ZN(n1411)
         );
  XNOR2_X1 U1531 ( .A(n287), .B(n1693), .ZN(n1278) );
  OAI22_X1 U1532 ( .A1(n1697), .A2(n1278), .B1(n307), .B2(n1277), .ZN(n1410)
         );
  XNOR2_X1 U1533 ( .A(n1279), .B(n1280), .ZN(n1282) );
  XNOR2_X1 U1534 ( .A(n1282), .B(n1281), .ZN(n1443) );
  FA_X1 U1535 ( .A(n1285), .B(n1284), .CI(n1283), .CO(n1301), .S(n1294) );
  FA_X1 U1536 ( .A(n1288), .B(n1287), .CI(n1286), .CO(n1293), .S(n1479) );
  XNOR2_X1 U1537 ( .A(n1294), .B(n1293), .ZN(n1289) );
  XNOR2_X1 U1538 ( .A(n1292), .B(n1289), .ZN(n1469) );
  OAI21_X1 U1539 ( .B1(n1467), .B2(n1468), .A(n1469), .ZN(n1291) );
  NOR2_X1 U1540 ( .A1(n1293), .A2(n1294), .ZN(n1297) );
  INV_X1 U1541 ( .A(n1292), .ZN(n1296) );
  NAND2_X1 U1542 ( .A1(n1294), .A2(n1293), .ZN(n1295) );
  OAI21_X1 U1543 ( .B1(n1297), .B2(n1296), .A(n1295), .ZN(n1348) );
  OR2_X1 U1544 ( .A1(n3555), .A2(n1901), .ZN(n1808) );
  NOR2_X1 U1545 ( .A1(n1809), .A2(n1808), .ZN(n1342) );
  FA_X1 U1546 ( .A(n1307), .B(n1306), .CI(n1305), .CO(n1562), .S(n1337) );
  XNOR2_X1 U1547 ( .A(xmem_data[31]), .B(fmem_data[4]), .ZN(n1501) );
  OAI22_X1 U1548 ( .A1(n234), .A2(n1308), .B1(n1501), .B2(n1743), .ZN(n1509)
         );
  XNOR2_X1 U1549 ( .A(n245), .B(n203), .ZN(n1494) );
  OAI22_X1 U1550 ( .A1(n196), .A2(n1309), .B1(n140), .B2(n1494), .ZN(n1508) );
  XNOR2_X1 U1551 ( .A(n258), .B(n1638), .ZN(n1500) );
  OR2_X1 U1552 ( .A1(n1500), .A2(n307), .ZN(n1310) );
  OAI21_X1 U1553 ( .B1(n1312), .B2(n1311), .A(n1310), .ZN(n1507) );
  FA_X1 U1554 ( .A(n1315), .B(n1314), .CI(n1313), .CO(n1505), .S(n1332) );
  XNOR2_X1 U1555 ( .A(fmem_data[6]), .B(n281), .ZN(n1493) );
  OAI22_X1 U1556 ( .A1(n1732), .A2(n1316), .B1(n1493), .B2(n1731), .ZN(n1542)
         );
  INV_X1 U1557 ( .A(n1542), .ZN(n1495) );
  XNOR2_X1 U1558 ( .A(fmem_data[14]), .B(n1530), .ZN(n1502) );
  OAI22_X1 U1559 ( .A1(n1585), .A2(n1317), .B1(n1584), .B2(n1502), .ZN(n1496)
         );
  XNOR2_X1 U1560 ( .A(n1495), .B(n1496), .ZN(n1320) );
  XNOR2_X1 U1561 ( .A(n1610), .B(fmem_data[12]), .ZN(n1510) );
  OR2_X1 U1562 ( .A1(n1510), .A2(n1641), .ZN(n1318) );
  OAI21_X1 U1563 ( .B1(n1008), .B2(n1319), .A(n1318), .ZN(n1497) );
  XNOR2_X1 U1564 ( .A(n1320), .B(n1497), .ZN(n1504) );
  FA_X1 U1565 ( .A(n1321), .B(n1323), .CI(n239), .CO(n1517), .S(n1329) );
  OAI22_X1 U1566 ( .A1(n1511), .A2(n1253), .B1(n199), .B2(n1325), .ZN(n1516)
         );
  FA_X1 U1567 ( .A(n1328), .B(n1327), .CI(n1326), .CO(n1515), .S(n1334) );
  FA_X1 U1568 ( .A(n1331), .B(n1330), .CI(n1329), .CO(n1491), .S(n1307) );
  OAI21_X1 U1569 ( .B1(n1334), .B2(n1333), .A(n1332), .ZN(n1336) );
  NAND2_X1 U1570 ( .A1(n1334), .A2(n200), .ZN(n1335) );
  NAND2_X1 U1571 ( .A1(n1336), .A2(n1335), .ZN(n1490) );
  XNOR2_X1 U1572 ( .A(n1946), .B(n1945), .ZN(n1810) );
  NOR2_X1 U1573 ( .A1(n1342), .A2(n299), .ZN(n1817) );
  XNOR2_X1 U1574 ( .A(n1901), .B(n3555), .ZN(n1805) );
  FA_X1 U1575 ( .A(n1345), .B(n1344), .CI(n1343), .CO(n1900), .S(n1959) );
  NOR2_X1 U1576 ( .A1(n1805), .A2(n1959), .ZN(n1807) );
  FA_X1 U1577 ( .A(n1348), .B(n1347), .CI(n1346), .CO(n1901), .S(n3556) );
  NOR2_X1 U1578 ( .A1(n3556), .A2(n187), .ZN(n1902) );
  NOR2_X1 U1579 ( .A1(n1807), .A2(n1902), .ZN(n1349) );
  NAND2_X1 U1580 ( .A1(n1817), .A2(n1349), .ZN(n1819) );
  FA_X1 U1581 ( .A(n1352), .B(n1350), .CI(n1351), .CO(n1258), .S(n1448) );
  OAI22_X1 U1582 ( .A1(n1356), .A2(n1355), .B1(n1354), .B2(n1353), .ZN(n1381)
         );
  OAI22_X1 U1583 ( .A1(n1008), .A2(n1358), .B1(n1357), .B2(n1641), .ZN(n1380)
         );
  OAI22_X1 U1584 ( .A1(n723), .A2(n1360), .B1(n141), .B2(n1359), .ZN(n1379) );
  XNOR2_X1 U1585 ( .A(n1362), .B(n1361), .ZN(n1364) );
  XNOR2_X1 U1586 ( .A(n1364), .B(n1363), .ZN(n1446) );
  FA_X1 U1587 ( .A(n1367), .B(n1366), .CI(n1365), .CO(n1442), .S(n1438) );
  XNOR2_X1 U1588 ( .A(n1369), .B(n1368), .ZN(n1409) );
  OAI22_X1 U1589 ( .A1(n1372), .A2(n1010), .B1(n297), .B2(n1370), .ZN(n1408)
         );
  FA_X1 U1590 ( .A(n1373), .B(n1374), .CI(n1375), .CO(n1407), .S(n1403) );
  INV_X1 U1591 ( .A(n1433), .ZN(n1384) );
  FA_X1 U1592 ( .A(n1378), .B(n1377), .CI(n1376), .CO(n1431), .S(n1426) );
  FA_X1 U1593 ( .A(n1381), .B(n1380), .CI(n1379), .CO(n1447), .S(n1430) );
  NOR2_X1 U1594 ( .A1(n1431), .A2(n1430), .ZN(n1383) );
  FA_X1 U1595 ( .A(n1387), .B(n1386), .CI(n1385), .CO(n1422), .S(n1464) );
  NAND2_X1 U1596 ( .A1(n1388), .A2(n1390), .ZN(n1393) );
  NAND2_X1 U1597 ( .A1(n1388), .A2(n1389), .ZN(n1392) );
  NAND2_X1 U1598 ( .A1(n1390), .A2(n1389), .ZN(n1391) );
  NAND3_X1 U1599 ( .A1(n1393), .A2(n1392), .A3(n1391), .ZN(n1415) );
  FA_X1 U1600 ( .A(n1396), .B(n1395), .CI(n1394), .CO(n1414), .S(n1401) );
  FA_X1 U1601 ( .A(n1399), .B(n1398), .CI(n1397), .CO(n1365), .S(n1413) );
  XNOR2_X1 U1602 ( .A(n1400), .B(n1413), .ZN(n1421) );
  FA_X1 U1603 ( .A(n1401), .B(n1402), .CI(n1403), .CO(n1420), .S(n1427) );
  OAI21_X2 U1604 ( .B1(n1406), .B2(n1405), .A(n1404), .ZN(n1455) );
  FA_X1 U1605 ( .A(n1409), .B(n1408), .CI(n1407), .CO(n1451), .S(n1433) );
  FA_X1 U1606 ( .A(n1412), .B(n1411), .CI(n1410), .CO(n1444), .S(n1450) );
  NAND2_X1 U1607 ( .A1(n1415), .A2(n1413), .ZN(n1418) );
  NAND2_X1 U1608 ( .A1(n1413), .A2(n1414), .ZN(n1417) );
  NAND2_X1 U1609 ( .A1(n1415), .A2(n1414), .ZN(n1416) );
  NAND3_X1 U1610 ( .A1(n1418), .A2(n1417), .A3(n1416), .ZN(n1449) );
  XNOR2_X1 U1611 ( .A(n1455), .B(n1454), .ZN(n1419) );
  XNOR2_X1 U1612 ( .A(n1453), .B(n1419), .ZN(n1799) );
  XNOR2_X1 U1613 ( .A(n1421), .B(n1420), .ZN(n1423) );
  XNOR2_X1 U1614 ( .A(n1423), .B(n1422), .ZN(n1461) );
  OR2_X1 U1615 ( .A1(n1427), .A2(n1426), .ZN(n1425) );
  NAND2_X1 U1616 ( .A1(n1425), .A2(n1424), .ZN(n1429) );
  NAND2_X1 U1617 ( .A1(n1427), .A2(n1426), .ZN(n1428) );
  NAND2_X1 U1618 ( .A1(n1429), .A2(n1428), .ZN(n1460) );
  NAND2_X1 U1619 ( .A1(n1461), .A2(n1460), .ZN(n1436) );
  XNOR2_X1 U1620 ( .A(n1433), .B(n1432), .ZN(n1459) );
  NAND2_X1 U1621 ( .A1(n1461), .A2(n1459), .ZN(n1435) );
  NAND2_X1 U1622 ( .A1(n1460), .A2(n1459), .ZN(n1434) );
  NAND3_X1 U1623 ( .A1(n1436), .A2(n1435), .A3(n1434), .ZN(n1798) );
  FA_X1 U1624 ( .A(n1439), .B(n1438), .CI(n1437), .CO(n1485), .S(n1453) );
  FA_X1 U1625 ( .A(n1442), .B(n1441), .CI(n1440), .CO(n1477), .S(n1484) );
  XNOR2_X1 U1626 ( .A(n1485), .B(n1484), .ZN(n1452) );
  FA_X1 U1627 ( .A(n1445), .B(n1444), .CI(n1443), .CO(n1474), .S(n1473) );
  FA_X1 U1628 ( .A(n1448), .B(n1447), .CI(n1446), .CO(n1472), .S(n1439) );
  FA_X1 U1629 ( .A(n1451), .B(n1450), .CI(n1449), .CO(n1471), .S(n1454) );
  XNOR2_X1 U1630 ( .A(n1452), .B(n1483), .ZN(n1801) );
  NAND2_X1 U1631 ( .A1(n1453), .A2(n1455), .ZN(n1458) );
  NAND2_X1 U1632 ( .A1(n1453), .A2(n1454), .ZN(n1457) );
  NAND2_X1 U1633 ( .A1(n1455), .A2(n1454), .ZN(n1456) );
  NAND3_X1 U1634 ( .A1(n1458), .A2(n1457), .A3(n1456), .ZN(n1800) );
  NAND2_X1 U1635 ( .A1(n2047), .A2(n2051), .ZN(n2026) );
  XOR2_X1 U1636 ( .A(n1460), .B(n1459), .Z(n1462) );
  XNOR2_X1 U1637 ( .A(n1462), .B(n1461), .ZN(n1795) );
  FA_X1 U1638 ( .A(n1465), .B(n1464), .CI(n1463), .CO(n1796), .S(n1087) );
  INV_X1 U1639 ( .A(n1796), .ZN(n1466) );
  NAND2_X1 U1640 ( .A1(n1795), .A2(n1466), .ZN(n2173) );
  INV_X1 U1641 ( .A(n2173), .ZN(n2030) );
  NOR2_X1 U1642 ( .A1(n2063), .A2(n2030), .ZN(n1488) );
  XNOR2_X1 U1643 ( .A(n1468), .B(n1467), .ZN(n1470) );
  XNOR2_X1 U1644 ( .A(n1470), .B(n1469), .ZN(n1876) );
  FA_X1 U1645 ( .A(n1473), .B(n1472), .CI(n1471), .CO(n1482), .S(n1483) );
  FA_X1 U1646 ( .A(n1476), .B(n1475), .CI(n1474), .CO(n1292), .S(n1481) );
  FA_X1 U1647 ( .A(n1479), .B(n1478), .CI(n1477), .CO(n1468), .S(n1480) );
  NOR2_X1 U1648 ( .A1(n1876), .A2(n1875), .ZN(n1803) );
  NAND2_X1 U1649 ( .A1(n1483), .A2(n341), .ZN(n1487) );
  NAND2_X1 U1650 ( .A1(n1485), .A2(n1484), .ZN(n1486) );
  NOR2_X1 U1651 ( .A1(n1878), .A2(n1877), .ZN(n2068) );
  NOR2_X1 U1652 ( .A1(n1803), .A2(n2068), .ZN(n3549) );
  NAND2_X1 U1653 ( .A1(n1488), .A2(n3549), .ZN(n1489) );
  NOR2_X1 U1654 ( .A1(n1819), .A2(n1489), .ZN(n1751) );
  FA_X1 U1655 ( .A(n1492), .B(n1491), .CI(n1490), .CO(n1559), .S(n1560) );
  XNOR2_X1 U1656 ( .A(fmem_data[7]), .B(n281), .ZN(n1528) );
  OAI22_X1 U1657 ( .A1(n1713), .A2(n1493), .B1(n1528), .B2(n1731), .ZN(n1543)
         );
  XNOR2_X1 U1658 ( .A(fmem_data[11]), .B(n246), .ZN(n1544) );
  OAI22_X1 U1659 ( .A1(n276), .A2(n1494), .B1(n140), .B2(n1544), .ZN(n1541) );
  OAI21_X1 U1660 ( .B1(n1497), .B2(n1496), .A(n1495), .ZN(n1499) );
  NAND2_X1 U1661 ( .A1(n1497), .A2(n1496), .ZN(n1498) );
  NAND2_X1 U1662 ( .A1(n1499), .A2(n1498), .ZN(n1520) );
  XNOR2_X1 U1663 ( .A(n184), .B(n1693), .ZN(n1549) );
  OAI22_X1 U1664 ( .A1(n1697), .A2(n1500), .B1(n307), .B2(n1549), .ZN(n1536)
         );
  XNOR2_X1 U1665 ( .A(xmem_data[31]), .B(fmem_data[5]), .ZN(n1546) );
  OAI22_X1 U1666 ( .A1(n234), .A2(n1501), .B1(n1546), .B2(n1743), .ZN(n1538)
         );
  XNOR2_X1 U1667 ( .A(fmem_data[15]), .B(n1530), .ZN(n1531) );
  OAI22_X1 U1668 ( .A1(n1585), .A2(n1502), .B1(n1533), .B2(n1531), .ZN(n1537)
         );
  XNOR2_X1 U1669 ( .A(n1538), .B(n1537), .ZN(n1503) );
  XNOR2_X1 U1670 ( .A(n1536), .B(n1503), .ZN(n1519) );
  FA_X1 U1671 ( .A(n1506), .B(n1505), .CI(n1504), .CO(n1551), .S(n1561) );
  FA_X1 U1672 ( .A(n1509), .B(n1508), .CI(n1507), .CO(n1523), .S(n1506) );
  XNOR2_X1 U1673 ( .A(n1610), .B(n194), .ZN(n1529) );
  OAI22_X1 U1674 ( .A1(n1008), .A2(n1510), .B1(n1529), .B2(n1641), .ZN(n1525)
         );
  AOI21_X1 U1675 ( .B1(n199), .B2(n1253), .A(n1511), .ZN(n1513) );
  INV_X1 U1676 ( .A(n1513), .ZN(n1524) );
  FA_X1 U1677 ( .A(n1517), .B(n1516), .CI(n1515), .CO(n1552), .S(n1492) );
  XNOR2_X1 U1678 ( .A(n1553), .B(n1552), .ZN(n1518) );
  XNOR2_X1 U1679 ( .A(n1551), .B(n1518), .ZN(n1557) );
  FA_X1 U1680 ( .A(n1521), .B(n1520), .CI(n1519), .CO(n1595), .S(n1558) );
  OR2_X1 U1681 ( .A1(n1525), .A2(n1524), .ZN(n1522) );
  NAND2_X1 U1682 ( .A1(n1523), .A2(n1522), .ZN(n1527) );
  NAND2_X1 U1683 ( .A1(n1525), .A2(n1524), .ZN(n1526) );
  NAND2_X1 U1684 ( .A1(n1527), .A2(n1526), .ZN(n1592) );
  XNOR2_X1 U1685 ( .A(fmem_data[8]), .B(n1711), .ZN(n1574) );
  OAI22_X1 U1686 ( .A1(n1732), .A2(n1528), .B1(n1574), .B2(n1731), .ZN(n1614)
         );
  INV_X1 U1687 ( .A(n1614), .ZN(n1589) );
  XNOR2_X1 U1688 ( .A(n1610), .B(fmem_data[14]), .ZN(n1573) );
  OAI22_X1 U1689 ( .A1(n1008), .A2(n1529), .B1(n1573), .B2(n1641), .ZN(n1588)
         );
  XNOR2_X1 U1690 ( .A(fmem_data[31]), .B(n1530), .ZN(n1583) );
  OAI22_X1 U1691 ( .A1(n1583), .A2(n1533), .B1(n1585), .B2(n1531), .ZN(n1587)
         );
  FA_X1 U1692 ( .A(n1543), .B(n1542), .CI(n1541), .CO(n1568), .S(n1521) );
  XNOR2_X1 U1693 ( .A(fmem_data[12]), .B(n182), .ZN(n1576) );
  OAI22_X1 U1694 ( .A1(n196), .A2(n1544), .B1(n140), .B2(n1576), .ZN(n1580) );
  XNOR2_X1 U1695 ( .A(xmem_data[31]), .B(fmem_data[6]), .ZN(n1572) );
  OR2_X1 U1696 ( .A1(n1572), .A2(n1743), .ZN(n1545) );
  OAI21_X1 U1697 ( .B1(n235), .B2(n1546), .A(n1545), .ZN(n1579) );
  XNOR2_X1 U1698 ( .A(n1579), .B(n1580), .ZN(n1550) );
  XNOR2_X1 U1699 ( .A(n203), .B(n1693), .ZN(n1570) );
  OR2_X1 U1700 ( .A1(n1570), .A2(n306), .ZN(n1548) );
  OAI21_X1 U1701 ( .B1(n1697), .B2(n1549), .A(n1548), .ZN(n1578) );
  XNOR2_X1 U1702 ( .A(n1550), .B(n1578), .ZN(n1567) );
  XNOR2_X1 U1703 ( .A(n1563), .B(n1564), .ZN(n1908) );
  XNOR2_X1 U1704 ( .A(n1908), .B(n1907), .ZN(n1975) );
  XNOR2_X1 U1705 ( .A(n1949), .B(n1975), .ZN(n1755) );
  FA_X1 U1706 ( .A(n1559), .B(n1558), .CI(n1557), .CO(n1949), .S(n1948) );
  FA_X1 U1707 ( .A(n1562), .B(n1561), .CI(n1560), .CO(n1947), .S(n1946) );
  OR2_X1 U1708 ( .A1(n1948), .A2(n1947), .ZN(n1754) );
  NOR2_X1 U1709 ( .A1(n1755), .A2(n1754), .ZN(n1598) );
  FA_X1 U1710 ( .A(n1569), .B(n1568), .CI(n1567), .CO(n1619), .S(n1564) );
  XNOR2_X1 U1711 ( .A(fmem_data[11]), .B(n1693), .ZN(n1605) );
  OAI22_X1 U1712 ( .A1(n1697), .A2(n1570), .B1(n306), .B2(n1605), .ZN(n1602)
         );
  BUF_X2 U1713 ( .A(n1571), .Z(n1747) );
  XNOR2_X1 U1714 ( .A(xmem_data[31]), .B(n238), .ZN(n1603) );
  OAI22_X1 U1715 ( .A1(n1747), .A2(n1572), .B1(n1603), .B2(n1743), .ZN(n1601)
         );
  XNOR2_X1 U1716 ( .A(n1610), .B(fmem_data[15]), .ZN(n1611) );
  OAI22_X1 U1717 ( .A1(n1008), .A2(n1573), .B1(n1611), .B2(n1641), .ZN(n1600)
         );
  XNOR2_X1 U1718 ( .A(fmem_data[9]), .B(n1711), .ZN(n1612) );
  OAI22_X1 U1719 ( .A1(n1732), .A2(n1574), .B1(n1731), .B2(n1612), .ZN(n1615)
         );
  XNOR2_X1 U1720 ( .A(n246), .B(fmem_data[13]), .ZN(n1604) );
  OAI22_X1 U1721 ( .A1(n274), .A2(n1576), .B1(n140), .B2(n1604), .ZN(n1613) );
  XNOR2_X1 U1722 ( .A(n1621), .B(n1620), .ZN(n1577) );
  XNOR2_X1 U1723 ( .A(n1619), .B(n1577), .ZN(n1624) );
  OAI21_X1 U1724 ( .B1(n1580), .B2(n1579), .A(n1578), .ZN(n1582) );
  NAND2_X1 U1725 ( .A1(n1579), .A2(n1580), .ZN(n1581) );
  AOI21_X1 U1726 ( .B1(n1585), .B2(n1584), .A(n1583), .ZN(n1586) );
  INV_X1 U1727 ( .A(n1586), .ZN(n1607) );
  FA_X1 U1728 ( .A(n1589), .B(n1588), .CI(n1587), .CO(n1606), .S(n1593) );
  XNOR2_X1 U1729 ( .A(n1624), .B(n1625), .ZN(n1597) );
  INV_X1 U1730 ( .A(n1593), .ZN(n1591) );
  INV_X1 U1731 ( .A(n1592), .ZN(n1590) );
  NAND2_X1 U1732 ( .A1(n1591), .A2(n1590), .ZN(n1594) );
  AOI22_X1 U1733 ( .A1(n1595), .A2(n1594), .B1(n1593), .B2(n1592), .ZN(n1596)
         );
  INV_X1 U1734 ( .A(n1596), .ZN(n1626) );
  XNOR2_X1 U1735 ( .A(n1597), .B(n1626), .ZN(n1910) );
  XNOR2_X1 U1736 ( .A(n1909), .B(n1910), .ZN(n1757) );
  OR2_X1 U1737 ( .A1(n1975), .A2(n1949), .ZN(n1756) );
  NOR2_X1 U1738 ( .A1(n1757), .A2(n1756), .ZN(n1760) );
  NOR2_X1 U1739 ( .A1(n1598), .A2(n1760), .ZN(n1763) );
  OR2_X1 U1740 ( .A1(n1945), .A2(n1946), .ZN(n1753) );
  XNOR2_X1 U1741 ( .A(n265), .B(n255), .ZN(n1752) );
  NAND2_X1 U1742 ( .A1(n1763), .A2(n1599), .ZN(n1750) );
  OR2_X1 U1743 ( .A1(n1910), .A2(n1909), .ZN(n1765) );
  FA_X1 U1744 ( .A(n1602), .B(n1601), .CI(n1600), .CO(n1635), .S(n1621) );
  XNOR2_X1 U1745 ( .A(xmem_data[31]), .B(n258), .ZN(n1640) );
  OAI22_X1 U1746 ( .A1(n1747), .A2(n1603), .B1(n1640), .B2(n1743), .ZN(n1649)
         );
  XNOR2_X1 U1747 ( .A(fmem_data[14]), .B(n182), .ZN(n1646) );
  OAI22_X1 U1748 ( .A1(n274), .A2(n1604), .B1(n191), .B2(n1646), .ZN(n1648) );
  XNOR2_X1 U1749 ( .A(fmem_data[12]), .B(n1693), .ZN(n1639) );
  OAI22_X1 U1750 ( .A1(n1697), .A2(n1605), .B1(n307), .B2(n1639), .ZN(n1647)
         );
  XNOR2_X1 U1751 ( .A(n1635), .B(n1634), .ZN(n1609) );
  FA_X1 U1752 ( .A(n1608), .B(n1607), .CI(n1606), .CO(n1633), .S(n1625) );
  XNOR2_X1 U1753 ( .A(n1609), .B(n1633), .ZN(n1655) );
  XNOR2_X1 U1754 ( .A(fmem_data[31]), .B(n1610), .ZN(n1642) );
  OAI22_X1 U1755 ( .A1(n1642), .A2(n1641), .B1(n1008), .B2(n1611), .ZN(n1652)
         );
  XNOR2_X1 U1756 ( .A(n203), .B(n1711), .ZN(n1645) );
  OAI22_X1 U1757 ( .A1(n1713), .A2(n1612), .B1(n1645), .B2(n1731), .ZN(n1663)
         );
  INV_X1 U1758 ( .A(n1663), .ZN(n1651) );
  FA_X1 U1759 ( .A(n1615), .B(n1613), .CI(n1614), .CO(n1650), .S(n1620) );
  INV_X1 U1760 ( .A(n1621), .ZN(n1617) );
  INV_X1 U1761 ( .A(n1620), .ZN(n1616) );
  NAND2_X1 U1762 ( .A1(n1617), .A2(n1616), .ZN(n1618) );
  NAND2_X1 U1763 ( .A1(n1619), .A2(n1618), .ZN(n1623) );
  NAND2_X1 U1764 ( .A1(n1623), .A2(n1622), .ZN(n1653) );
  BUF_X1 U1765 ( .A(n1937), .Z(n1629) );
  XNOR2_X1 U1766 ( .A(n1629), .B(n1938), .ZN(n1764) );
  NOR2_X1 U1767 ( .A1(n1765), .A2(n1764), .ZN(n1673) );
  OR2_X1 U1768 ( .A1(n1629), .A2(n1938), .ZN(n1767) );
  INV_X1 U1769 ( .A(n1635), .ZN(n1631) );
  INV_X1 U1770 ( .A(n1634), .ZN(n1630) );
  NAND2_X1 U1771 ( .A1(n1631), .A2(n1630), .ZN(n1632) );
  NAND2_X1 U1772 ( .A1(n1633), .A2(n1632), .ZN(n1637) );
  NAND2_X1 U1773 ( .A1(n1635), .A2(n1634), .ZN(n1636) );
  NAND2_X1 U1774 ( .A1(n1637), .A2(n1636), .ZN(n1671) );
  XNOR2_X1 U1775 ( .A(n194), .B(n1693), .ZN(n1659) );
  OAI22_X1 U1776 ( .A1(n1697), .A2(n1639), .B1(n306), .B2(n1659), .ZN(n1668)
         );
  XNOR2_X1 U1777 ( .A(xmem_data[31]), .B(n184), .ZN(n1660) );
  OAI22_X1 U1778 ( .A1(n1747), .A2(n1640), .B1(n1660), .B2(n1743), .ZN(n1667)
         );
  NAND2_X1 U1779 ( .A1(n1008), .A2(n1641), .ZN(n1644) );
  INV_X1 U1780 ( .A(n1642), .ZN(n1643) );
  NAND2_X1 U1781 ( .A1(n1644), .A2(n1643), .ZN(n1666) );
  XNOR2_X1 U1782 ( .A(fmem_data[11]), .B(n1711), .ZN(n1661) );
  OAI22_X1 U1783 ( .A1(n1713), .A2(n1645), .B1(n1661), .B2(n1731), .ZN(n1664)
         );
  XNOR2_X1 U1784 ( .A(fmem_data[15]), .B(n246), .ZN(n1665) );
  OAI22_X1 U1785 ( .A1(n276), .A2(n1646), .B1(n191), .B2(n1665), .ZN(n1662) );
  FA_X1 U1786 ( .A(n1649), .B(n1648), .CI(n1647), .CO(n1657), .S(n1634) );
  FA_X1 U1787 ( .A(n1652), .B(n1651), .CI(n1650), .CO(n1656), .S(n1654) );
  FA_X1 U1788 ( .A(n1655), .B(n1654), .CI(n1653), .CO(n1939), .S(n1937) );
  XNOR2_X1 U1789 ( .A(n216), .B(n1939), .ZN(n1766) );
  OR2_X1 U1790 ( .A1(n1767), .A2(n1766), .ZN(n1672) );
  OR2_X1 U1791 ( .A1(n216), .A2(n1939), .ZN(n1769) );
  XNOR2_X1 U1792 ( .A(n188), .B(n1693), .ZN(n1682) );
  OAI22_X1 U1793 ( .A1(n1697), .A2(n1659), .B1(n307), .B2(n1682), .ZN(n1685)
         );
  XNOR2_X1 U1794 ( .A(xmem_data[31]), .B(n203), .ZN(n1678) );
  OAI22_X1 U1795 ( .A1(n234), .A2(n1660), .B1(n1678), .B2(n1743), .ZN(n1684)
         );
  XNOR2_X1 U1796 ( .A(fmem_data[12]), .B(n281), .ZN(n1677) );
  OAI22_X1 U1797 ( .A1(n1713), .A2(n1661), .B1(n1677), .B2(n1731), .ZN(n1705)
         );
  INV_X1 U1798 ( .A(n1705), .ZN(n1683) );
  FA_X1 U1799 ( .A(n1664), .B(n1663), .CI(n1662), .CO(n1676), .S(n1658) );
  XNOR2_X1 U1800 ( .A(fmem_data[31]), .B(n195), .ZN(n1679) );
  OAI22_X1 U1801 ( .A1(n1679), .A2(n191), .B1(n196), .B2(n1665), .ZN(n1675) );
  FA_X1 U1802 ( .A(n1668), .B(n1667), .CI(n1666), .CO(n1674), .S(n1670) );
  FA_X1 U1803 ( .A(n1671), .B(n1670), .CI(n1669), .CO(n1941), .S(n1940) );
  XNOR2_X1 U1804 ( .A(n278), .B(n137), .ZN(n1768) );
  NAND2_X1 U1805 ( .A1(n1672), .A2(n1771), .ZN(n1775) );
  NOR2_X1 U1806 ( .A1(n1673), .A2(n1775), .ZN(n1745) );
  OR2_X1 U1807 ( .A1(n278), .A2(n137), .ZN(n1777) );
  FA_X1 U1808 ( .A(n1676), .B(n1675), .CI(n1674), .CO(n1725), .S(n1686) );
  XNOR2_X1 U1809 ( .A(n194), .B(n281), .ZN(n1691) );
  OAI22_X1 U1810 ( .A1(n1713), .A2(n1677), .B1(n1691), .B2(n256), .ZN(n1706)
         );
  XNOR2_X1 U1811 ( .A(xmem_data[31]), .B(fmem_data[11]), .ZN(n1692) );
  OAI22_X1 U1812 ( .A1(n234), .A2(n1678), .B1(n1692), .B2(n1743), .ZN(n1704)
         );
  AOI21_X1 U1813 ( .B1(n274), .B2(n140), .A(n1679), .ZN(n1681) );
  INV_X1 U1814 ( .A(n1681), .ZN(n1709) );
  XNOR2_X1 U1815 ( .A(n192), .B(n1693), .ZN(n1694) );
  OAI22_X1 U1816 ( .A1(n1697), .A2(n1682), .B1(n306), .B2(n1694), .ZN(n1708)
         );
  FA_X1 U1817 ( .A(n1685), .B(n1684), .CI(n1683), .CO(n1707), .S(n1687) );
  FA_X1 U1818 ( .A(n1688), .B(n1687), .CI(n1686), .CO(n2001), .S(n1942) );
  XNOR2_X1 U1819 ( .A(n2002), .B(n2001), .ZN(n1776) );
  NOR2_X1 U1820 ( .A1(n1777), .A2(n1776), .ZN(n1690) );
  NOR2_X1 U1821 ( .A1(n1690), .A2(n1689), .ZN(n1738) );
  XNOR2_X1 U1822 ( .A(n188), .B(n281), .ZN(n1699) );
  OAI22_X1 U1823 ( .A1(n1713), .A2(n1691), .B1(n1699), .B2(n1731), .ZN(n1715)
         );
  INV_X1 U1824 ( .A(n1715), .ZN(n1703) );
  XNOR2_X1 U1825 ( .A(xmem_data[31]), .B(fmem_data[12]), .ZN(n1700) );
  OAI22_X1 U1826 ( .A1(n235), .A2(n1692), .B1(n1700), .B2(n1743), .ZN(n1702)
         );
  XNOR2_X1 U1827 ( .A(fmem_data[31]), .B(n1693), .ZN(n1695) );
  OAI22_X1 U1828 ( .A1(n1695), .A2(n306), .B1(n1697), .B2(n1694), .ZN(n1701)
         );
  AOI21_X1 U1829 ( .B1(n1697), .B2(n307), .A(n1695), .ZN(n1698) );
  INV_X1 U1830 ( .A(n1698), .ZN(n1718) );
  XNOR2_X1 U1831 ( .A(fmem_data[15]), .B(n1711), .ZN(n1712) );
  OAI22_X1 U1832 ( .A1(n1713), .A2(n1699), .B1(n1712), .B2(n256), .ZN(n1716)
         );
  XNOR2_X1 U1833 ( .A(xmem_data[31]), .B(n194), .ZN(n1710) );
  OAI22_X1 U1834 ( .A1(n1747), .A2(n1700), .B1(n1710), .B2(n1743), .ZN(n1714)
         );
  FA_X1 U1835 ( .A(n1703), .B(n1702), .CI(n1701), .CO(n1719), .S(n1722) );
  FA_X1 U1836 ( .A(n1706), .B(n1705), .CI(n1704), .CO(n1721), .S(n1724) );
  FA_X1 U1837 ( .A(n1709), .B(n1708), .CI(n1707), .CO(n1720), .S(n1723) );
  XNOR2_X1 U1838 ( .A(xmem_data[31]), .B(n188), .ZN(n1729) );
  OAI22_X1 U1839 ( .A1(n235), .A2(n1710), .B1(n1729), .B2(n1743), .ZN(n1740)
         );
  INV_X1 U1840 ( .A(n1740), .ZN(n1736) );
  XNOR2_X1 U1841 ( .A(fmem_data[31]), .B(n281), .ZN(n1730) );
  OAI22_X1 U1842 ( .A1(n1730), .A2(n256), .B1(n1713), .B2(n1712), .ZN(n1735)
         );
  FA_X1 U1843 ( .A(n1716), .B(n1715), .CI(n1714), .CO(n1734), .S(n1717) );
  FA_X1 U1844 ( .A(n1719), .B(n1718), .CI(n1717), .CO(n1916), .S(n1915) );
  NOR2_X1 U1845 ( .A1(n340), .A2(n308), .ZN(n1781) );
  FA_X1 U1846 ( .A(n1722), .B(n1721), .CI(n1720), .CO(n1914), .S(n1913) );
  INV_X1 U1847 ( .A(n1913), .ZN(n1727) );
  FA_X1 U1848 ( .A(n1725), .B(n1724), .CI(n1723), .CO(n1912), .S(n2002) );
  INV_X1 U1849 ( .A(n1912), .ZN(n1726) );
  NAND2_X1 U1850 ( .A1(n1727), .A2(n1726), .ZN(n1728) );
  NAND2_X1 U1851 ( .A1(n1781), .A2(n1728), .ZN(n1737) );
  XNOR2_X1 U1852 ( .A(xmem_data[31]), .B(n192), .ZN(n1742) );
  OAI22_X1 U1853 ( .A1(n1747), .A2(n1729), .B1(n1742), .B2(n231), .ZN(n1741)
         );
  AOI21_X1 U1854 ( .B1(n1713), .B2(n256), .A(n1730), .ZN(n1733) );
  INV_X1 U1855 ( .A(n1733), .ZN(n1739) );
  FA_X1 U1856 ( .A(n1736), .B(n1735), .CI(n1734), .CO(n1919), .S(n1917) );
  NOR2_X1 U1857 ( .A1(n1737), .A2(n310), .ZN(n1784) );
  NAND2_X1 U1858 ( .A1(n1738), .A2(n1784), .ZN(n1744) );
  FA_X1 U1859 ( .A(n1741), .B(n1740), .CI(n1739), .CO(n1927), .S(n1920) );
  XNOR2_X1 U1860 ( .A(fmem_data[31]), .B(xmem_data[31]), .ZN(n1746) );
  OAI22_X1 U1861 ( .A1(n1746), .A2(n1743), .B1(n234), .B2(n1742), .ZN(n1929)
         );
  INV_X1 U1862 ( .A(n1929), .ZN(n1926) );
  NOR2_X1 U1863 ( .A1(n1744), .A2(n311), .ZN(n1788) );
  NAND2_X1 U1864 ( .A1(n1745), .A2(n1788), .ZN(n1791) );
  AOI21_X1 U1865 ( .B1(n235), .B2(n231), .A(n1746), .ZN(n1748) );
  INV_X1 U1866 ( .A(n1748), .ZN(n1930) );
  OR2_X1 U1867 ( .A1(n1930), .A2(n1929), .ZN(n1793) );
  NAND2_X1 U1868 ( .A1(n1751), .A2(n1821), .ZN(n1825) );
  AND2_X1 U1869 ( .A1(n1753), .A2(n1752), .ZN(n1762) );
  NAND2_X1 U1870 ( .A1(n1755), .A2(n1754), .ZN(n1759) );
  NAND2_X1 U1871 ( .A1(n1757), .A2(n1756), .ZN(n1758) );
  OAI21_X1 U1872 ( .B1(n1760), .B2(n1759), .A(n1758), .ZN(n1761) );
  AOI21_X1 U1873 ( .B1(n1763), .B2(n1762), .A(n1761), .ZN(n1792) );
  NAND2_X1 U1874 ( .A1(n1765), .A2(n1764), .ZN(n1774) );
  AND2_X1 U1875 ( .A1(n1767), .A2(n1766), .ZN(n1772) );
  AND2_X1 U1876 ( .A1(n1769), .A2(n1768), .ZN(n1770) );
  AOI21_X1 U1877 ( .B1(n1772), .B2(n1771), .A(n1770), .ZN(n1773) );
  OAI21_X1 U1878 ( .B1(n1775), .B2(n1774), .A(n1773), .ZN(n1789) );
  NAND2_X1 U1879 ( .A1(n1777), .A2(n1776), .ZN(n1778) );
  OAI21_X1 U1880 ( .B1(n1778), .B2(n1689), .A(n335), .ZN(n1785) );
  XNOR2_X1 U1881 ( .A(n1915), .B(n1914), .ZN(n1780) );
  OAI21_X1 U1882 ( .B1(n337), .B2(n308), .A(n314), .ZN(n1779) );
  AOI21_X1 U1883 ( .B1(n1781), .B2(n1780), .A(n1779), .ZN(n1782) );
  OAI21_X1 U1884 ( .B1(n1782), .B2(n310), .A(n338), .ZN(n1783) );
  AOI21_X1 U1885 ( .B1(n1785), .B2(n1784), .A(n1783), .ZN(n1786) );
  OAI21_X1 U1886 ( .B1(n1786), .B2(n311), .A(n332), .ZN(n1787) );
  AOI21_X1 U1887 ( .B1(n1789), .B2(n1788), .A(n1787), .ZN(n1790) );
  OAI21_X1 U1888 ( .B1(n1792), .B2(n1791), .A(n1790), .ZN(n1794) );
  NAND2_X1 U1889 ( .A1(n1794), .A2(n1793), .ZN(n1824) );
  INV_X1 U1890 ( .A(n1795), .ZN(n1797) );
  NAND2_X1 U1891 ( .A1(n1797), .A2(n1796), .ZN(n2172) );
  NAND2_X1 U1892 ( .A1(n1799), .A2(n1798), .ZN(n2058) );
  INV_X1 U1893 ( .A(n2058), .ZN(n2048) );
  AND2_X1 U1894 ( .A1(n1801), .A2(n1800), .ZN(n2034) );
  AOI21_X1 U1895 ( .B1(n2051), .B2(n2048), .A(n2034), .ZN(n1802) );
  OAI21_X1 U1896 ( .B1(n2063), .B2(n2172), .A(n1802), .ZN(n1804) );
  NAND2_X1 U1897 ( .A1(n1878), .A2(n1877), .ZN(n2069) );
  NAND2_X1 U1898 ( .A1(n1876), .A2(n1875), .ZN(n2041) );
  OAI21_X1 U1899 ( .B1(n1803), .B2(n2069), .A(n2041), .ZN(n3547) );
  AOI21_X1 U1900 ( .B1(n1804), .B2(n3549), .A(n3547), .ZN(n1820) );
  NAND2_X1 U1901 ( .A1(n3556), .A2(n187), .ZN(n1962) );
  NAND2_X1 U1902 ( .A1(n1805), .A2(n1959), .ZN(n1806) );
  OAI21_X1 U1903 ( .B1(n1807), .B2(n1962), .A(n1806), .ZN(n1816) );
  NAND2_X1 U1904 ( .A1(n1809), .A2(n1808), .ZN(n1813) );
  NAND2_X1 U1905 ( .A1(n1811), .A2(n1810), .ZN(n1812) );
  OAI21_X1 U1906 ( .B1(n1814), .B2(n1813), .A(n1812), .ZN(n1815) );
  AOI21_X1 U1907 ( .B1(n251), .B2(n1816), .A(n1815), .ZN(n1818) );
  OAI21_X1 U1908 ( .B1(n1820), .B2(n1819), .A(n1818), .ZN(n1822) );
  NAND2_X1 U1909 ( .A1(n1822), .A2(n254), .ZN(n1823) );
  NAND2_X1 U1910 ( .A1(\ctrl_conv_output_inst/conv_start_accum ), .A2(n4009), 
        .ZN(n1827) );
  NAND2_X1 U1911 ( .A1(conv_pre_start), .A2(n4102), .ZN(n2604) );
  INV_X1 U1912 ( .A(n2604), .ZN(n4010) );
  NAND2_X1 U1913 ( .A1(n3291), .A2(n4010), .ZN(n2022) );
  INV_X1 U1914 ( .A(n2022), .ZN(n3562) );
  NAND2_X1 U1915 ( .A1(n3561), .A2(n3562), .ZN(n2025) );
  BUF_X2 U1916 ( .A(n2025), .Z(n2203) );
  INV_X1 U1917 ( .A(n2093), .ZN(n1842) );
  INV_X1 U1918 ( .A(n237), .ZN(n2158) );
  NOR2_X1 U1919 ( .A1(n2164), .A2(n3651), .ZN(n1838) );
  INV_X1 U1920 ( .A(n1830), .ZN(n2114) );
  INV_X1 U1921 ( .A(n1831), .ZN(n2197) );
  INV_X1 U1922 ( .A(n1832), .ZN(n2198) );
  INV_X1 U1923 ( .A(n2196), .ZN(n1833) );
  AOI21_X1 U1924 ( .B1(n2197), .B2(n2198), .A(n1833), .ZN(n2221) );
  OAI21_X1 U1925 ( .B1(n1834), .B2(n2221), .A(n2219), .ZN(n2115) );
  INV_X1 U1926 ( .A(n2113), .ZN(n1835) );
  AOI21_X1 U1927 ( .B1(n2114), .B2(n2115), .A(n1835), .ZN(n2109) );
  OAI21_X1 U1928 ( .B1(n2109), .B2(n1836), .A(n2106), .ZN(n3650) );
  OAI21_X1 U1929 ( .B1(n2164), .B2(n3652), .A(n2165), .ZN(n1837) );
  OAI21_X1 U1930 ( .B1(n2183), .B2(n2179), .A(n2180), .ZN(n2081) );
  INV_X1 U1931 ( .A(n2084), .ZN(n1839) );
  NOR2_X1 U1932 ( .A1(n2082), .A2(n1839), .ZN(n1841) );
  OAI21_X1 U1933 ( .B1(n1839), .B2(n2099), .A(n2083), .ZN(n1840) );
  AOI21_X1 U1934 ( .B1(n2081), .B2(n1841), .A(n1840), .ZN(n2090) );
  OAI21_X1 U1935 ( .B1(n1842), .B2(n3645), .A(n2092), .ZN(n2155) );
  INV_X1 U1936 ( .A(n2157), .ZN(n1843) );
  AOI21_X1 U1937 ( .B1(n2155), .B2(n2158), .A(n1843), .ZN(n1844) );
  OAI21_X1 U1938 ( .B1(n1845), .B2(n2090), .A(n1844), .ZN(n2120) );
  INV_X1 U1939 ( .A(n1846), .ZN(n2141) );
  INV_X1 U1940 ( .A(n2139), .ZN(n3641) );
  NAND2_X1 U1941 ( .A1(n2141), .A2(n3641), .ZN(n2122) );
  NOR2_X1 U1942 ( .A1(n1849), .A2(n2122), .ZN(n1851) );
  INV_X1 U1943 ( .A(n3640), .ZN(n1848) );
  INV_X1 U1944 ( .A(n2140), .ZN(n1847) );
  AOI21_X1 U1945 ( .B1(n2141), .B2(n1848), .A(n1847), .ZN(n2121) );
  OAI21_X1 U1946 ( .B1(n2121), .B2(n1849), .A(n2123), .ZN(n1850) );
  AOI21_X1 U1947 ( .B1(n2120), .B2(n1851), .A(n1850), .ZN(n2147) );
  INV_X1 U1948 ( .A(n2133), .ZN(n1853) );
  INV_X1 U1949 ( .A(n2075), .ZN(n2130) );
  NOR2_X1 U1950 ( .A1(n1853), .A2(n2130), .ZN(n1856) );
  NAND2_X1 U1951 ( .A1(n1856), .A2(n1852), .ZN(n1858) );
  AOI21_X1 U1952 ( .B1(n1856), .B2(n1855), .A(n1854), .ZN(n1857) );
  OAI21_X1 U1953 ( .B1(n1879), .B2(n3670), .A(n3663), .ZN(n2032) );
  INV_X1 U1954 ( .A(n2032), .ZN(n1860) );
  NAND2_X1 U1955 ( .A1(n1874), .A2(n185), .ZN(n1862) );
  XNOR2_X1 U1956 ( .A(n1863), .B(n1862), .ZN(n2023) );
  NAND2_X1 U1957 ( .A1(n2149), .A2(n236), .ZN(n1867) );
  NOR2_X1 U1958 ( .A1(n1867), .A2(n1869), .ZN(n1873) );
  AOI21_X1 U1959 ( .B1(n2149), .B2(n263), .A(n211), .ZN(n1870) );
  OAI21_X1 U1960 ( .B1(n1870), .B2(n1869), .A(n298), .ZN(n1871) );
  AOI21_X1 U1961 ( .B1(n1872), .B2(n1873), .A(n1871), .ZN(n1898) );
  NAND2_X1 U1962 ( .A1(n1874), .A2(n2173), .ZN(n1891) );
  INV_X1 U1963 ( .A(n1891), .ZN(n1881) );
  NAND2_X1 U1964 ( .A1(n2047), .A2(n2051), .ZN(n2063) );
  NOR2_X1 U1965 ( .A1(n1885), .A2(n2026), .ZN(n1893) );
  INV_X1 U1966 ( .A(n1879), .ZN(n3664) );
  INV_X1 U1967 ( .A(n3660), .ZN(n3671) );
  AND2_X1 U1968 ( .A1(n3664), .A2(n3671), .ZN(n1880) );
  NAND3_X1 U1969 ( .A1(n1893), .A2(n1881), .A3(n1880), .ZN(n1897) );
  AOI21_X1 U1970 ( .B1(n2051), .B2(n2048), .A(n2034), .ZN(n1884) );
  INV_X1 U1971 ( .A(n2069), .ZN(n1882) );
  NAND2_X1 U1972 ( .A1(n1882), .A2(n2042), .ZN(n1883) );
  OAI211_X1 U1973 ( .C1(n1885), .C2(n1884), .A(n2041), .B(n1883), .ZN(n1886)
         );
  INV_X1 U1974 ( .A(n1886), .ZN(n1896) );
  INV_X1 U1975 ( .A(n3670), .ZN(n1888) );
  INV_X1 U1976 ( .A(n3663), .ZN(n1887) );
  AOI21_X1 U1977 ( .B1(n3664), .B2(n1888), .A(n1887), .ZN(n1892) );
  INV_X1 U1978 ( .A(n2029), .ZN(n1889) );
  AOI21_X1 U1979 ( .B1(n1889), .B2(n2173), .A(n293), .ZN(n1890) );
  OAI21_X1 U1980 ( .B1(n1892), .B2(n1891), .A(n1890), .ZN(n1894) );
  NAND2_X1 U1981 ( .A1(n1894), .A2(n222), .ZN(n1895) );
  OAI211_X1 U1982 ( .C1(n1898), .C2(n1897), .A(n1896), .B(n1895), .ZN(n2021)
         );
  AND2_X1 U1983 ( .A1(n1901), .A2(n3555), .ZN(n1964) );
  NOR2_X1 U1984 ( .A1(n1965), .A2(n1964), .ZN(n1958) );
  INV_X1 U1985 ( .A(n1945), .ZN(n1899) );
  XNOR2_X1 U1986 ( .A(n1946), .B(n1899), .ZN(n1967) );
  AND2_X1 U1987 ( .A1(n288), .A2(n1900), .ZN(n1966) );
  NOR2_X1 U1988 ( .A1(n1967), .A2(n1966), .ZN(n1957) );
  NOR2_X1 U1989 ( .A1(n1957), .A2(n1958), .ZN(n1905) );
  XNOR2_X1 U1990 ( .A(n187), .B(n1901), .ZN(n1960) );
  NOR2_X1 U1991 ( .A1(n1960), .A2(n1959), .ZN(n1903) );
  NOR2_X1 U1992 ( .A1(n1903), .A2(n1902), .ZN(n1904) );
  NAND2_X1 U1993 ( .A1(n1905), .A2(n1904), .ZN(n1956) );
  INV_X1 U1994 ( .A(n1909), .ZN(n1906) );
  XNOR2_X1 U1995 ( .A(n1910), .B(n1906), .ZN(n1982) );
  XNOR2_X1 U1996 ( .A(n1908), .B(n1907), .ZN(n1950) );
  AND2_X1 U1997 ( .A1(n1950), .A2(n1949), .ZN(n1981) );
  OR2_X1 U1998 ( .A1(n1982), .A2(n1981), .ZN(n1911) );
  NAND2_X1 U1999 ( .A1(n1911), .A2(n1986), .ZN(n1989) );
  INV_X1 U2000 ( .A(n1989), .ZN(n1955) );
  HA_X1 U2001 ( .A(n1913), .B(n1912), .S(n2003) );
  INV_X1 U2002 ( .A(n2003), .ZN(n2006) );
  HA_X1 U2003 ( .A(n1915), .B(n1914), .S(n1925) );
  HA_X1 U2004 ( .A(n1917), .B(n1916), .S(n1918) );
  INV_X1 U2005 ( .A(n1918), .ZN(n1923) );
  HA_X1 U2006 ( .A(n1920), .B(n1919), .S(n1921) );
  INV_X1 U2007 ( .A(n1921), .ZN(n1922) );
  NOR2_X1 U2008 ( .A1(n1923), .A2(n1922), .ZN(n1924) );
  NAND2_X1 U2009 ( .A1(n1925), .A2(n1924), .ZN(n1935) );
  HA_X1 U2010 ( .A(n1927), .B(n1926), .S(n1928) );
  INV_X1 U2011 ( .A(n1928), .ZN(n1933) );
  HA_X1 U2012 ( .A(n1930), .B(n1929), .S(n1931) );
  INV_X1 U2013 ( .A(n1931), .ZN(n1932) );
  OR2_X1 U2014 ( .A1(n1933), .A2(n1932), .ZN(n1934) );
  NOR2_X1 U2015 ( .A1(n1935), .A2(n1934), .ZN(n2009) );
  NAND2_X1 U2016 ( .A1(n1936), .A2(n2009), .ZN(n2011) );
  HA_X1 U2017 ( .A(n1937), .B(n1938), .CO(n1992), .S(n1984) );
  OR2_X1 U2018 ( .A1(n1993), .A2(n1992), .ZN(n1943) );
  HA_X1 U2019 ( .A(n1940), .B(n1939), .CO(n1995), .S(n1993) );
  HA_X1 U2020 ( .A(n1942), .B(n1941), .CO(n2000), .S(n1994) );
  NAND2_X1 U2021 ( .A1(n1943), .A2(n1997), .ZN(n1991) );
  NOR2_X1 U2022 ( .A1(n2011), .A2(n1991), .ZN(n1954) );
  INV_X1 U2023 ( .A(n1947), .ZN(n1944) );
  XNOR2_X1 U2024 ( .A(n1944), .B(n1948), .ZN(n1973) );
  OR2_X1 U2025 ( .A1(n1973), .A2(n334), .ZN(n1953) );
  INV_X1 U2026 ( .A(n1976), .ZN(n1952) );
  INV_X1 U2027 ( .A(n1949), .ZN(n1974) );
  NAND2_X1 U2028 ( .A1(n1952), .A2(n1951), .ZN(n1978) );
  NOR2_X1 U2029 ( .A1(n1956), .A2(n2017), .ZN(n2020) );
  NOR2_X1 U2030 ( .A1(n1960), .A2(n1959), .ZN(n1963) );
  NAND2_X1 U2031 ( .A1(n1960), .A2(n1959), .ZN(n1961) );
  OAI21_X1 U2032 ( .B1(n1963), .B2(n1962), .A(n1961), .ZN(n1972) );
  INV_X1 U2033 ( .A(n1967), .ZN(n1970) );
  NAND2_X1 U2034 ( .A1(n1965), .A2(n1964), .ZN(n1969) );
  NAND2_X1 U2035 ( .A1(n1967), .A2(n1966), .ZN(n1968) );
  OAI21_X1 U2036 ( .B1(n1970), .B2(n1969), .A(n1968), .ZN(n1971) );
  AOI21_X1 U2037 ( .B1(n1972), .B2(n1905), .A(n1971), .ZN(n2018) );
  AND2_X1 U2038 ( .A1(n334), .A2(n1973), .ZN(n1980) );
  XNOR2_X1 U2039 ( .A(n1975), .B(n1974), .ZN(n1977) );
  AND2_X1 U2040 ( .A1(n1976), .A2(n1977), .ZN(n1979) );
  OAI21_X1 U2041 ( .B1(n1980), .B2(n1979), .A(n1978), .ZN(n1990) );
  AND2_X1 U2042 ( .A1(n1982), .A2(n1981), .ZN(n1987) );
  AND2_X1 U2043 ( .A1(n1984), .A2(n1983), .ZN(n1985) );
  AOI21_X1 U2044 ( .B1(n1987), .B2(n1986), .A(n1985), .ZN(n1988) );
  OAI21_X1 U2045 ( .B1(n1990), .B2(n1989), .A(n1988), .ZN(n2015) );
  NOR2_X1 U2046 ( .A1(n2011), .A2(n1991), .ZN(n2014) );
  AND2_X1 U2047 ( .A1(n1993), .A2(n1992), .ZN(n1998) );
  AND2_X1 U2048 ( .A1(n1995), .A2(n1994), .ZN(n1996) );
  AOI21_X1 U2049 ( .B1(n1997), .B2(n1998), .A(n1996), .ZN(n2012) );
  NAND2_X1 U2050 ( .A1(n2000), .A2(n1999), .ZN(n2007) );
  HA_X1 U2051 ( .A(n2002), .B(n2001), .CO(n2004), .S(n1999) );
  NAND2_X1 U2052 ( .A1(n2004), .A2(n2003), .ZN(n2005) );
  OAI21_X1 U2053 ( .B1(n2007), .B2(n2006), .A(n2005), .ZN(n2008) );
  NAND2_X1 U2054 ( .A1(n2009), .A2(n2008), .ZN(n2010) );
  OAI21_X1 U2055 ( .B1(n2012), .B2(n2011), .A(n2010), .ZN(n2013) );
  AOI21_X1 U2056 ( .B1(n2015), .B2(n2014), .A(n2013), .ZN(n2016) );
  OAI21_X1 U2057 ( .B1(n2018), .B2(n2017), .A(n2016), .ZN(n2019) );
  AOI21_X1 U2058 ( .B1(n2021), .B2(n2020), .A(n2019), .ZN(n3565) );
  NOR2_X1 U2059 ( .A1(n3565), .A2(n2022), .ZN(n2055) );
  BUF_X2 U2060 ( .A(n2055), .Z(n3657) );
  NAND2_X1 U2061 ( .A1(n2023), .A2(n3668), .ZN(n2024) );
  NAND3_X1 U2062 ( .A1(n2203), .A2(n2024), .A3(n342), .ZN(\mac_unit_inst/n138 ) );
  INV_X1 U2063 ( .A(n3661), .ZN(n3673) );
  NOR2_X1 U2064 ( .A1(n2063), .A2(n2068), .ZN(n2038) );
  NOR2_X1 U2065 ( .A1(n2030), .A2(n2027), .ZN(n2033) );
  NAND2_X1 U2066 ( .A1(n2028), .A2(n2033), .ZN(n3546) );
  INV_X1 U2067 ( .A(n3546), .ZN(n2064) );
  NAND2_X1 U2068 ( .A1(n2038), .A2(n2064), .ZN(n2040) );
  OAI21_X1 U2069 ( .B1(n2030), .B2(n185), .A(n2172), .ZN(n2031) );
  INV_X1 U2070 ( .A(n3552), .ZN(n2065) );
  NAND2_X1 U2071 ( .A1(n2048), .A2(n2051), .ZN(n2035) );
  INV_X1 U2072 ( .A(n2034), .ZN(n2052) );
  NAND2_X1 U2073 ( .A1(n2035), .A2(n2052), .ZN(n3548) );
  INV_X1 U2074 ( .A(n3548), .ZN(n2036) );
  OAI21_X1 U2075 ( .B1(n2036), .B2(n2068), .A(n268), .ZN(n2037) );
  AOI21_X1 U2076 ( .B1(n2065), .B2(n2038), .A(n2037), .ZN(n2039) );
  OAI21_X1 U2077 ( .B1(n3673), .B2(n2040), .A(n2039), .ZN(n2044) );
  NAND2_X1 U2078 ( .A1(n2042), .A2(n2041), .ZN(n2043) );
  XNOR2_X1 U2079 ( .A(n2044), .B(n2043), .ZN(n2045) );
  BUF_X2 U2080 ( .A(n2055), .Z(n3668) );
  NAND2_X1 U2081 ( .A1(n2045), .A2(n3680), .ZN(n2046) );
  NAND3_X1 U2082 ( .A1(n3681), .A2(n2046), .A3(n343), .ZN(\mac_unit_inst/n143 ) );
  NAND2_X1 U2083 ( .A1(n292), .A2(n3562), .ZN(n2074) );
  BUF_X2 U2084 ( .A(n2074), .Z(n3658) );
  NAND2_X1 U2085 ( .A1(n2064), .A2(n2047), .ZN(n2050) );
  AOI21_X1 U2086 ( .B1(n2065), .B2(n2047), .A(n2048), .ZN(n2049) );
  OAI21_X1 U2087 ( .B1(n3673), .B2(n2050), .A(n2049), .ZN(n2054) );
  NAND2_X1 U2088 ( .A1(n2051), .A2(n2052), .ZN(n2053) );
  XNOR2_X1 U2089 ( .A(n2054), .B(n2053), .ZN(n2056) );
  BUF_X2 U2090 ( .A(n2055), .Z(n3680) );
  NAND2_X1 U2091 ( .A1(n2056), .A2(n3668), .ZN(n2057) );
  NAND3_X1 U2092 ( .A1(n3658), .A2(n2057), .A3(n344), .ZN(\mac_unit_inst/n141 ) );
  OAI21_X1 U2093 ( .B1(n3673), .B2(n3546), .A(n3552), .ZN(n2060) );
  NAND2_X1 U2094 ( .A1(n2047), .A2(n2058), .ZN(n2059) );
  XNOR2_X1 U2095 ( .A(n2060), .B(n2059), .ZN(n2061) );
  NAND2_X1 U2096 ( .A1(n2061), .A2(n3668), .ZN(n2062) );
  NAND3_X1 U2097 ( .A1(n2062), .A2(n3658), .A3(n345), .ZN(\mac_unit_inst/n140 ) );
  INV_X1 U2098 ( .A(n2063), .ZN(n3545) );
  NAND2_X1 U2099 ( .A1(n2064), .A2(n3545), .ZN(n2067) );
  AOI21_X1 U2100 ( .B1(n2065), .B2(n3545), .A(n3548), .ZN(n2066) );
  OAI21_X1 U2101 ( .B1(n3673), .B2(n2067), .A(n2066), .ZN(n2071) );
  NAND2_X1 U2102 ( .A1(n301), .A2(n268), .ZN(n2070) );
  XNOR2_X1 U2103 ( .A(n2071), .B(n2070), .ZN(n2072) );
  BUF_X2 U2104 ( .A(n2074), .Z(n2227) );
  NAND2_X1 U2105 ( .A1(n2075), .A2(n139), .ZN(n2077) );
  XOR2_X1 U2106 ( .A(n218), .B(n2077), .Z(n2079) );
  NOR2_X1 U2107 ( .A1(n2223), .A2(n4141), .ZN(n2078) );
  AOI21_X1 U2108 ( .B1(n3680), .B2(n2079), .A(n2078), .ZN(n2080) );
  NAND2_X1 U2109 ( .A1(n2227), .A2(n2080), .ZN(\mac_unit_inst/n134 ) );
  INV_X1 U2110 ( .A(n2081), .ZN(n2102) );
  OAI21_X1 U2111 ( .B1(n2102), .B2(n2082), .A(n2099), .ZN(n2086) );
  NAND2_X1 U2112 ( .A1(n2084), .A2(n2083), .ZN(n2085) );
  XNOR2_X1 U2113 ( .A(n2086), .B(n2085), .ZN(n2088) );
  NOR2_X1 U2114 ( .A1(n3659), .A2(n4126), .ZN(n2087) );
  INV_X1 U2115 ( .A(n186), .ZN(n3648) );
  AOI21_X1 U2116 ( .B1(n3648), .B2(n3646), .A(n2091), .ZN(n2095) );
  NAND2_X1 U2117 ( .A1(n2093), .A2(n2092), .ZN(n2094) );
  XOR2_X1 U2118 ( .A(n2095), .B(n2094), .Z(n2097) );
  NOR2_X1 U2119 ( .A1(n3659), .A2(n4124), .ZN(n2096) );
  NAND2_X1 U2120 ( .A1(n2100), .A2(n2099), .ZN(n2101) );
  XOR2_X1 U2121 ( .A(n2102), .B(n2101), .Z(n2104) );
  NOR2_X1 U2122 ( .A1(n3659), .A2(n4127), .ZN(n2103) );
  NAND2_X1 U2123 ( .A1(n2107), .A2(n2106), .ZN(n2108) );
  XOR2_X1 U2124 ( .A(n2109), .B(n2108), .Z(n2111) );
  NOR2_X1 U2125 ( .A1(n3659), .A2(n4131), .ZN(n2110) );
  AOI21_X1 U2126 ( .B1(n3680), .B2(n2111), .A(n2110), .ZN(n2112) );
  NAND2_X1 U2127 ( .A1(n2227), .A2(n2112), .ZN(\mac_unit_inst/n120 ) );
  NAND2_X1 U2128 ( .A1(n2114), .A2(n2113), .ZN(n2116) );
  XNOR2_X1 U2129 ( .A(n2116), .B(n2115), .ZN(n2118) );
  NOR2_X1 U2130 ( .A1(n3659), .A2(n4114), .ZN(n2117) );
  AOI21_X1 U2131 ( .B1(n3668), .B2(n2118), .A(n2117), .ZN(n2119) );
  NAND2_X1 U2132 ( .A1(n2227), .A2(n2119), .ZN(\mac_unit_inst/n119 ) );
  INV_X1 U2133 ( .A(n2120), .ZN(n3643) );
  OAI21_X1 U2134 ( .B1(n3643), .B2(n2122), .A(n2121), .ZN(n2126) );
  NAND2_X1 U2135 ( .A1(n2124), .A2(n2123), .ZN(n2125) );
  XNOR2_X1 U2136 ( .A(n2126), .B(n2125), .ZN(n2128) );
  NOR2_X1 U2137 ( .A1(n3659), .A2(n4120), .ZN(n2127) );
  AOI21_X1 U2138 ( .B1(n3668), .B2(n2128), .A(n2127), .ZN(n2129) );
  NAND2_X1 U2139 ( .A1(n2227), .A2(n2129), .ZN(\mac_unit_inst/n131 ) );
  OAI21_X1 U2140 ( .B1(n218), .B2(n2130), .A(n139), .ZN(n2135) );
  NAND2_X1 U2141 ( .A1(n2133), .A2(n2132), .ZN(n2134) );
  XNOR2_X1 U2142 ( .A(n2135), .B(n2134), .ZN(n2137) );
  NOR2_X1 U2143 ( .A1(n2223), .A2(n4140), .ZN(n2136) );
  OAI21_X1 U2144 ( .B1(n3643), .B2(n2139), .A(n294), .ZN(n2143) );
  NAND2_X1 U2145 ( .A1(n2141), .A2(n2140), .ZN(n2142) );
  XNOR2_X1 U2146 ( .A(n2143), .B(n2142), .ZN(n2145) );
  NOR2_X1 U2147 ( .A1(n3659), .A2(n4121), .ZN(n2144) );
  AOI21_X1 U2148 ( .B1(n3668), .B2(n2145), .A(n2144), .ZN(n2146) );
  NAND2_X1 U2149 ( .A1(n2203), .A2(n2146), .ZN(\mac_unit_inst/n130 ) );
  INV_X1 U2150 ( .A(n303), .ZN(n3678) );
  AOI21_X1 U2151 ( .B1(n3678), .B2(n236), .A(n263), .ZN(n2151) );
  NAND2_X1 U2152 ( .A1(n2149), .A2(n2148), .ZN(n2150) );
  XOR2_X1 U2153 ( .A(n2151), .B(n2150), .Z(n2153) );
  NOR2_X1 U2154 ( .A1(n2223), .A2(n4142), .ZN(n2152) );
  AOI21_X1 U2155 ( .B1(n3668), .B2(n2153), .A(n2152), .ZN(n2154) );
  NAND2_X1 U2156 ( .A1(n2203), .A2(n2154), .ZN(\mac_unit_inst/n133 ) );
  AOI21_X1 U2157 ( .B1(n3648), .B2(n2156), .A(n2155), .ZN(n2160) );
  NAND2_X1 U2158 ( .A1(n2158), .A2(n2157), .ZN(n2159) );
  XOR2_X1 U2159 ( .A(n2160), .B(n2159), .Z(n2162) );
  NOR2_X1 U2160 ( .A1(n3659), .A2(n4123), .ZN(n2161) );
  INV_X1 U2161 ( .A(n2164), .ZN(n2166) );
  NAND2_X1 U2162 ( .A1(n2166), .A2(n2165), .ZN(n2167) );
  XNOR2_X1 U2163 ( .A(n2168), .B(n2167), .ZN(n2170) );
  NOR2_X1 U2164 ( .A1(n3659), .A2(n4129), .ZN(n2169) );
  NAND2_X1 U2165 ( .A1(n2173), .A2(n2172), .ZN(n2174) );
  XNOR2_X1 U2166 ( .A(n2175), .B(n2174), .ZN(n2177) );
  NOR2_X1 U2167 ( .A1(n2223), .A2(n4136), .ZN(n2176) );
  AOI21_X1 U2168 ( .B1(n3680), .B2(n2177), .A(n2176), .ZN(n2178) );
  NAND2_X1 U2169 ( .A1(n2227), .A2(n2178), .ZN(\mac_unit_inst/n139 ) );
  INV_X1 U2170 ( .A(n2179), .ZN(n2181) );
  NAND2_X1 U2171 ( .A1(n2181), .A2(n2180), .ZN(n2182) );
  XOR2_X1 U2172 ( .A(n2183), .B(n2182), .Z(n2185) );
  NOR2_X1 U2173 ( .A1(n3659), .A2(n4128), .ZN(n2184) );
  AOI21_X1 U2174 ( .B1(n3668), .B2(n2185), .A(n2184), .ZN(n2186) );
  NAND2_X1 U2175 ( .A1(n2227), .A2(n2186), .ZN(\mac_unit_inst/n123 ) );
  AND2_X1 U2176 ( .A1(n284), .A2(xmem_data[0]), .ZN(n2188) );
  NOR2_X1 U2177 ( .A1(n2223), .A2(n4144), .ZN(n2187) );
  AOI21_X1 U2178 ( .B1(n3668), .B2(n2188), .A(n2187), .ZN(n2189) );
  NAND2_X1 U2179 ( .A1(n2227), .A2(n2189), .ZN(\mac_unit_inst/n113 ) );
  OR2_X1 U2180 ( .A1(n2191), .A2(n2190), .ZN(n2192) );
  AND2_X1 U2181 ( .A1(n2192), .A2(n2207), .ZN(n2194) );
  NOR2_X1 U2182 ( .A1(n2223), .A2(n4119), .ZN(n2193) );
  NAND2_X1 U2183 ( .A1(n2197), .A2(n2196), .ZN(n2199) );
  XNOR2_X1 U2184 ( .A(n2199), .B(n2198), .ZN(n2201) );
  NOR2_X1 U2185 ( .A1(n2223), .A2(n4116), .ZN(n2200) );
  AOI21_X1 U2186 ( .B1(n3657), .B2(n2201), .A(n2200), .ZN(n2202) );
  NAND2_X1 U2187 ( .A1(n2203), .A2(n2202), .ZN(\mac_unit_inst/n117 ) );
  INV_X1 U2188 ( .A(n2204), .ZN(n2206) );
  NAND2_X1 U2189 ( .A1(n2206), .A2(n2205), .ZN(n2208) );
  XOR2_X1 U2190 ( .A(n2208), .B(n2207), .Z(n2210) );
  NOR2_X1 U2191 ( .A1(n2223), .A2(n4118), .ZN(n2209) );
  AOI21_X1 U2192 ( .B1(n3668), .B2(n2210), .A(n2209), .ZN(n2211) );
  NAND2_X1 U2193 ( .A1(n2227), .A2(n2211), .ZN(\mac_unit_inst/n115 ) );
  NAND2_X1 U2194 ( .A1(n2213), .A2(n2212), .ZN(n2215) );
  XNOR2_X1 U2195 ( .A(n2215), .B(n2214), .ZN(n2217) );
  NOR2_X1 U2196 ( .A1(n2223), .A2(n4117), .ZN(n2216) );
  AOI21_X1 U2197 ( .B1(n3680), .B2(n2217), .A(n2216), .ZN(n2218) );
  NAND2_X1 U2198 ( .A1(n2227), .A2(n2218), .ZN(\mac_unit_inst/n116 ) );
  NAND2_X1 U2199 ( .A1(n2220), .A2(n2219), .ZN(n2222) );
  XOR2_X1 U2200 ( .A(n2222), .B(n2221), .Z(n2225) );
  NOR2_X1 U2201 ( .A1(n2223), .A2(n4115), .ZN(n2224) );
  AOI21_X1 U2202 ( .B1(n3668), .B2(n2225), .A(n2224), .ZN(n2226) );
  NAND2_X1 U2203 ( .A1(n2227), .A2(n2226), .ZN(\mac_unit_inst/n118 ) );
  NAND2_X1 U2204 ( .A1(n3779), .A2(n4105), .ZN(n2261) );
  NOR2_X1 U2205 ( .A1(n4070), .A2(n4082), .ZN(n3722) );
  NAND2_X1 U2206 ( .A1(xmem_addr[3]), .A2(n3722), .ZN(n2253) );
  NOR2_X1 U2207 ( .A1(n2261), .A2(n2253), .ZN(n3250) );
  NAND2_X1 U2208 ( .A1(n4070), .A2(n4082), .ZN(n2237) );
  NAND2_X1 U2209 ( .A1(xmem_addr[3]), .A2(n3710), .ZN(n2251) );
  NOR2_X1 U2210 ( .A1(n2261), .A2(n2251), .ZN(n3586) );
  AOI22_X1 U2211 ( .A1(n3574), .A2(\xmem_inst/mem[27][20] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][20] ), .ZN(n2231) );
  NOR2_X1 U2212 ( .A1(n2263), .A2(n2253), .ZN(n3254) );
  NAND2_X1 U2213 ( .A1(xmem_addr[5]), .A2(xmem_addr[2]), .ZN(n2264) );
  NAND2_X1 U2214 ( .A1(n4070), .A2(xmem_addr[0]), .ZN(n2236) );
  NAND2_X1 U2215 ( .A1(n3714), .A2(n4083), .ZN(n2259) );
  NOR2_X1 U2216 ( .A1(n2264), .A2(n2259), .ZN(n3184) );
  AOI22_X1 U2217 ( .A1(n3624), .A2(\xmem_inst/mem[11][20] ), .B1(n3613), .B2(
        \xmem_inst/mem[37][20] ), .ZN(n2230) );
  NAND2_X1 U2218 ( .A1(n3722), .A2(n4083), .ZN(n2258) );
  NOR2_X1 U2219 ( .A1(n2258), .A2(n2267), .ZN(n2967) );
  NAND2_X1 U2220 ( .A1(xmem_addr[3]), .A2(n3714), .ZN(n2262) );
  NOR2_X1 U2221 ( .A1(n2261), .A2(n2262), .ZN(n3147) );
  AOI22_X1 U2222 ( .A1(n3614), .A2(\xmem_inst/mem[23][20] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][20] ), .ZN(n2229) );
  NAND2_X1 U2223 ( .A1(n3710), .A2(n4083), .ZN(n2265) );
  NOR2_X1 U2224 ( .A1(n2265), .A2(n2263), .ZN(n3598) );
  NOR2_X1 U2225 ( .A1(n2267), .A2(n2262), .ZN(n3573) );
  AOI22_X1 U2226 ( .A1(n3233), .A2(\xmem_inst/mem[0][20] ), .B1(n3244), .B2(
        \xmem_inst/mem[29][20] ), .ZN(n2228) );
  NAND4_X1 U2227 ( .A1(n2231), .A2(n2230), .A3(n2229), .A4(n2228), .ZN(n2250)
         );
  NOR2_X1 U2228 ( .A1(xmem_addr[0]), .A2(n4070), .ZN(n3718) );
  NAND2_X1 U2229 ( .A1(n3718), .A2(n4083), .ZN(n2243) );
  NOR2_X1 U2230 ( .A1(n2243), .A2(n2267), .ZN(n3581) );
  NAND2_X1 U2231 ( .A1(xmem_addr[3]), .A2(n3718), .ZN(n2266) );
  NOR2_X1 U2232 ( .A1(n2261), .A2(n2266), .ZN(n3208) );
  AOI22_X1 U2233 ( .A1(n3581), .A2(\xmem_inst/mem[22][20] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][20] ), .ZN(n2235) );
  NAND2_X1 U2234 ( .A1(xmem_addr[5]), .A2(n4105), .ZN(n2260) );
  NOR2_X1 U2235 ( .A1(n2260), .A2(n2243), .ZN(n2958) );
  NOR2_X1 U2236 ( .A1(n2243), .A2(n2263), .ZN(n3234) );
  AOI22_X1 U2237 ( .A1(n3631), .A2(\xmem_inst/mem[34][20] ), .B1(n3615), .B2(
        \xmem_inst/mem[2][20] ), .ZN(n2234) );
  NAND2_X1 U2238 ( .A1(xmem_addr[2]), .A2(n3728), .ZN(n2252) );
  NOR2_X1 U2239 ( .A1(n2252), .A2(n2253), .ZN(n3618) );
  NOR2_X1 U2240 ( .A1(n2243), .A2(n2261), .ZN(n3153) );
  AOI22_X1 U2241 ( .A1(n3252), .A2(\xmem_inst/mem[15][20] ), .B1(n3568), .B2(
        \xmem_inst/mem[18][20] ), .ZN(n2233) );
  NOR2_X1 U2242 ( .A1(n2252), .A2(n2259), .ZN(n3567) );
  NOR2_X1 U2243 ( .A1(n2252), .A2(n2262), .ZN(n3210) );
  AOI22_X1 U2244 ( .A1(n3225), .A2(\xmem_inst/mem[5][20] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][20] ), .ZN(n2232) );
  NAND4_X1 U2245 ( .A1(n2235), .A2(n2234), .A3(n2233), .A4(n2232), .ZN(n2249)
         );
  NOR2_X1 U2246 ( .A1(n2243), .A2(n2252), .ZN(n3235) );
  NAND2_X1 U2247 ( .A1(xmem_addr[3]), .A2(xmem_addr[5]), .ZN(n2240) );
  NOR2_X1 U2248 ( .A1(n2236), .A2(n2240), .ZN(n3592) );
  AOI22_X1 U2249 ( .A1(n3235), .A2(\xmem_inst/mem[6][20] ), .B1(n3190), .B2(
        \xmem_inst/mem[41][20] ), .ZN(n2239) );
  NOR2_X1 U2250 ( .A1(n2252), .A2(n2266), .ZN(n3154) );
  NOR2_X1 U2251 ( .A1(n2237), .A2(n2240), .ZN(n2972) );
  AOI22_X1 U2252 ( .A1(n3616), .A2(\xmem_inst/mem[14][20] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][20] ), .ZN(n2238) );
  NAND2_X1 U2253 ( .A1(n2239), .A2(n2238), .ZN(n2248) );
  NOR2_X1 U2254 ( .A1(n2260), .A2(n2265), .ZN(n3148) );
  OR2_X1 U2255 ( .A1(n2258), .A2(n2252), .ZN(n3082) );
  NOR2_X1 U2256 ( .A1(n4070), .A2(n2240), .ZN(n3617) );
  NAND2_X1 U2257 ( .A1(n3245), .A2(\xmem_inst/mem[42][20] ), .ZN(n2241) );
  OAI21_X1 U2258 ( .B1(n3082), .B2(n4106), .A(n2241), .ZN(n2242) );
  AOI21_X1 U2259 ( .B1(n3602), .B2(\xmem_inst/mem[32][20] ), .A(n2242), .ZN(
        n2246) );
  OR2_X1 U2260 ( .A1(n2258), .A2(n2264), .ZN(n3114) );
  INV_X2 U2261 ( .A(n3114), .ZN(n3627) );
  NOR2_X1 U2262 ( .A1(n2267), .A2(n2251), .ZN(n3189) );
  AOI22_X1 U2263 ( .A1(n3627), .A2(\xmem_inst/mem[39][20] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][20] ), .ZN(n2245) );
  NOR2_X1 U2264 ( .A1(n2264), .A2(n2243), .ZN(n3203) );
  AOI22_X1 U2265 ( .A1(n3580), .A2(\xmem_inst/mem[38][20] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][20] ), .ZN(n2244) );
  NAND3_X1 U2266 ( .A1(n2246), .A2(n2245), .A3(n2244), .ZN(n2247) );
  OR4_X1 U2267 ( .A1(n2250), .A2(n2249), .A3(n2248), .A4(n2247), .ZN(n2274) );
  NOR2_X1 U2268 ( .A1(n2263), .A2(n2251), .ZN(n3591) );
  NOR2_X1 U2269 ( .A1(n2252), .A2(n2251), .ZN(n3177) );
  AOI22_X1 U2270 ( .A1(n3179), .A2(\xmem_inst/mem[8][20] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][20] ), .ZN(n2257) );
  NOR2_X1 U2271 ( .A1(n2265), .A2(n2252), .ZN(n3202) );
  NOR2_X1 U2272 ( .A1(n2261), .A2(n2259), .ZN(n3209) );
  AOI22_X1 U2273 ( .A1(n3604), .A2(\xmem_inst/mem[4][20] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][20] ), .ZN(n2256) );
  NOR2_X4 U2274 ( .A1(n2267), .A2(n2259), .ZN(n3600) );
  NOR2_X1 U2275 ( .A1(n2263), .A2(n2259), .ZN(n2295) );
  AOI22_X1 U2276 ( .A1(n3600), .A2(\xmem_inst/mem[21][20] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][20] ), .ZN(n2255) );
  OR2_X1 U2277 ( .A1(n2258), .A2(n2260), .ZN(n3021) );
  INV_X2 U2278 ( .A(n3021), .ZN(n3597) );
  NOR2_X1 U2279 ( .A1(n2267), .A2(n2253), .ZN(n3072) );
  AOI22_X1 U2280 ( .A1(n3597), .A2(\xmem_inst/mem[35][20] ), .B1(n3072), .B2(
        \xmem_inst/mem[31][20] ), .ZN(n2254) );
  NAND4_X1 U2281 ( .A1(n2257), .A2(n2256), .A3(n2255), .A4(n2254), .ZN(n2273)
         );
  NOR2_X4 U2282 ( .A1(n2258), .A2(n2263), .ZN(n3626) );
  NOR2_X1 U2283 ( .A1(n2260), .A2(n2259), .ZN(n3599) );
  AOI22_X1 U2284 ( .A1(n3626), .A2(\xmem_inst/mem[3][20] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][20] ), .ZN(n2271) );
  NOR2_X1 U2285 ( .A1(n2265), .A2(n2261), .ZN(n3084) );
  NOR2_X1 U2286 ( .A1(n2263), .A2(n2266), .ZN(n3603) );
  AOI22_X1 U2287 ( .A1(n3084), .A2(\xmem_inst/mem[16][20] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][20] ), .ZN(n2270) );
  NOR2_X1 U2288 ( .A1(n2263), .A2(n2262), .ZN(n3219) );
  NOR2_X1 U2289 ( .A1(n2264), .A2(n2265), .ZN(n3579) );
  AOI22_X1 U2290 ( .A1(n3619), .A2(\xmem_inst/mem[9][20] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][20] ), .ZN(n2269) );
  NOR2_X1 U2291 ( .A1(n2265), .A2(n2267), .ZN(n3251) );
  NOR2_X1 U2292 ( .A1(n2267), .A2(n2266), .ZN(n3178) );
  AOI22_X1 U2293 ( .A1(n3584), .A2(\xmem_inst/mem[20][20] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][20] ), .ZN(n2268) );
  NAND4_X1 U2294 ( .A1(n2271), .A2(n2270), .A3(n2269), .A4(n2268), .ZN(n2272)
         );
  OR3_X1 U2295 ( .A1(n2274), .A2(n2273), .A3(n2272), .ZN(\xmem_inst/N259 ) );
  AOI22_X1 U2296 ( .A1(n3598), .A2(\xmem_inst/mem[0][7] ), .B1(n3584), .B2(
        \xmem_inst/mem[20][7] ), .ZN(n2278) );
  AOI22_X1 U2297 ( .A1(n3568), .A2(\xmem_inst/mem[18][7] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][7] ), .ZN(n2277) );
  AOI22_X1 U2298 ( .A1(n3574), .A2(\xmem_inst/mem[27][7] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][7] ), .ZN(n2276) );
  AOI22_X1 U2299 ( .A1(n3627), .A2(\xmem_inst/mem[39][7] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][7] ), .ZN(n2275) );
  NAND4_X1 U2300 ( .A1(n2278), .A2(n2277), .A3(n2276), .A4(n2275), .ZN(n2294)
         );
  AOI22_X1 U2301 ( .A1(n3252), .A2(\xmem_inst/mem[15][7] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][7] ), .ZN(n2282) );
  AOI22_X1 U2302 ( .A1(n3616), .A2(\xmem_inst/mem[14][7] ), .B1(n3220), .B2(
        \xmem_inst/mem[36][7] ), .ZN(n2281) );
  AOI22_X1 U2303 ( .A1(n3614), .A2(\xmem_inst/mem[23][7] ), .B1(n3615), .B2(
        \xmem_inst/mem[2][7] ), .ZN(n2280) );
  AOI22_X1 U2304 ( .A1(n3193), .A2(\xmem_inst/mem[22][7] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][7] ), .ZN(n2279) );
  NAND4_X1 U2305 ( .A1(n2282), .A2(n2281), .A3(n2280), .A4(n2279), .ZN(n2293)
         );
  AOI22_X1 U2306 ( .A1(n3235), .A2(\xmem_inst/mem[6][7] ), .B1(n3244), .B2(
        \xmem_inst/mem[29][7] ), .ZN(n2286) );
  AOI22_X1 U2307 ( .A1(n3631), .A2(\xmem_inst/mem[34][7] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][7] ), .ZN(n2285) );
  AOI22_X1 U2308 ( .A1(n3600), .A2(\xmem_inst/mem[21][7] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][7] ), .ZN(n2284) );
  AOI22_X1 U2309 ( .A1(n3626), .A2(\xmem_inst/mem[3][7] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][7] ), .ZN(n2283) );
  NAND4_X1 U2310 ( .A1(n2286), .A2(n2285), .A3(n2284), .A4(n2283), .ZN(n2292)
         );
  AOI22_X1 U2311 ( .A1(n3190), .A2(\xmem_inst/mem[41][7] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][7] ), .ZN(n2290) );
  NAND2_X1 U2312 ( .A1(n3245), .A2(\xmem_inst/mem[42][7] ), .ZN(n2289) );
  NAND2_X1 U2313 ( .A1(n3601), .A2(\xmem_inst/mem[26][7] ), .ZN(n2288) );
  NAND2_X1 U2314 ( .A1(n3179), .A2(\xmem_inst/mem[8][7] ), .ZN(n2287) );
  NAND4_X1 U2315 ( .A1(n2290), .A2(n2289), .A3(n2288), .A4(n2287), .ZN(n2291)
         );
  OR4_X1 U2316 ( .A1(n2294), .A2(n2293), .A3(n2292), .A4(n2291), .ZN(n2305) );
  AOI22_X1 U2317 ( .A1(n3148), .A2(\xmem_inst/mem[32][7] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][7] ), .ZN(n2299) );
  AOI22_X1 U2318 ( .A1(n3597), .A2(\xmem_inst/mem[35][7] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][7] ), .ZN(n2298) );
  AOI22_X1 U2319 ( .A1(n3613), .A2(\xmem_inst/mem[37][7] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][7] ), .ZN(n2297) );
  BUF_X1 U2320 ( .A(n2295), .Z(n3628) );
  AOI22_X1 U2321 ( .A1(n3254), .A2(\xmem_inst/mem[11][7] ), .B1(n3628), .B2(
        \xmem_inst/mem[1][7] ), .ZN(n2296) );
  NAND4_X1 U2322 ( .A1(n2299), .A2(n2298), .A3(n2297), .A4(n2296), .ZN(n2304)
         );
  AOI22_X1 U2323 ( .A1(n3594), .A2(\xmem_inst/mem[19][7] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][7] ), .ZN(n2302) );
  AOI22_X1 U2324 ( .A1(n3629), .A2(\xmem_inst/mem[31][7] ), .B1(n3593), .B2(
        \xmem_inst/mem[40][7] ), .ZN(n2301) );
  AOI22_X1 U2325 ( .A1(n3580), .A2(\xmem_inst/mem[38][7] ), .B1(n3084), .B2(
        \xmem_inst/mem[16][7] ), .ZN(n2300) );
  NAND3_X1 U2326 ( .A1(n2302), .A2(n2301), .A3(n2300), .ZN(n2303) );
  OR3_X1 U2327 ( .A1(n2305), .A2(n2304), .A3(n2303), .ZN(\xmem_inst/N272 ) );
  AOI22_X1 U2328 ( .A1(n3602), .A2(\xmem_inst/mem[32][14] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][14] ), .ZN(n2309) );
  AOI22_X1 U2329 ( .A1(n3627), .A2(\xmem_inst/mem[39][14] ), .B1(n3604), .B2(
        \xmem_inst/mem[4][14] ), .ZN(n2308) );
  AOI22_X1 U2330 ( .A1(n3570), .A2(\xmem_inst/mem[17][14] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][14] ), .ZN(n2307) );
  AOI22_X1 U2331 ( .A1(n3235), .A2(\xmem_inst/mem[6][14] ), .B1(n3584), .B2(
        \xmem_inst/mem[20][14] ), .ZN(n2306) );
  NAND4_X1 U2332 ( .A1(n2309), .A2(n2308), .A3(n2307), .A4(n2306), .ZN(n2325)
         );
  AOI22_X1 U2333 ( .A1(n3233), .A2(\xmem_inst/mem[0][14] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][14] ), .ZN(n2313) );
  AOI22_X1 U2334 ( .A1(n3614), .A2(\xmem_inst/mem[23][14] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][14] ), .ZN(n2312) );
  AOI22_X1 U2335 ( .A1(n3628), .A2(\xmem_inst/mem[1][14] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][14] ), .ZN(n2311) );
  AOI22_X1 U2336 ( .A1(n3615), .A2(\xmem_inst/mem[2][14] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][14] ), .ZN(n2310) );
  NAND4_X1 U2337 ( .A1(n2313), .A2(n2312), .A3(n2311), .A4(n2310), .ZN(n2324)
         );
  AOI22_X1 U2338 ( .A1(n3582), .A2(\xmem_inst/mem[7][14] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][14] ), .ZN(n2317) );
  AOI22_X1 U2339 ( .A1(n3096), .A2(\xmem_inst/mem[10][14] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][14] ), .ZN(n2316) );
  AOI22_X1 U2340 ( .A1(n3574), .A2(\xmem_inst/mem[27][14] ), .B1(n3252), .B2(
        \xmem_inst/mem[15][14] ), .ZN(n2315) );
  AOI22_X1 U2341 ( .A1(n3624), .A2(\xmem_inst/mem[11][14] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][14] ), .ZN(n2314) );
  NAND4_X1 U2342 ( .A1(n2317), .A2(n2316), .A3(n2315), .A4(n2314), .ZN(n2323)
         );
  AOI22_X1 U2343 ( .A1(n3631), .A2(\xmem_inst/mem[34][14] ), .B1(n3190), .B2(
        \xmem_inst/mem[41][14] ), .ZN(n2321) );
  NAND2_X1 U2344 ( .A1(n3245), .A2(\xmem_inst/mem[42][14] ), .ZN(n2320) );
  NAND2_X1 U2345 ( .A1(n3616), .A2(\xmem_inst/mem[14][14] ), .ZN(n2319) );
  NAND2_X1 U2346 ( .A1(n3220), .A2(\xmem_inst/mem[36][14] ), .ZN(n2318) );
  NAND4_X1 U2347 ( .A1(n2321), .A2(n2320), .A3(n2319), .A4(n2318), .ZN(n2322)
         );
  OR4_X1 U2348 ( .A1(n2325), .A2(n2324), .A3(n2323), .A4(n2322), .ZN(n2335) );
  AOI22_X1 U2349 ( .A1(n3629), .A2(\xmem_inst/mem[31][14] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][14] ), .ZN(n2329) );
  AOI22_X1 U2350 ( .A1(n3580), .A2(\xmem_inst/mem[38][14] ), .B1(n3244), .B2(
        \xmem_inst/mem[29][14] ), .ZN(n2328) );
  AOI22_X1 U2351 ( .A1(n3626), .A2(\xmem_inst/mem[3][14] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][14] ), .ZN(n2327) );
  AOI22_X1 U2352 ( .A1(n3568), .A2(\xmem_inst/mem[18][14] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][14] ), .ZN(n2326) );
  NAND4_X1 U2353 ( .A1(n2329), .A2(n2328), .A3(n2327), .A4(n2326), .ZN(n2334)
         );
  AOI22_X1 U2354 ( .A1(n3597), .A2(\xmem_inst/mem[35][14] ), .B1(n3572), .B2(
        \xmem_inst/mem[25][14] ), .ZN(n2332) );
  AOI22_X1 U2355 ( .A1(n3594), .A2(\xmem_inst/mem[19][14] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][14] ), .ZN(n2331) );
  AOI22_X1 U2356 ( .A1(n3613), .A2(\xmem_inst/mem[37][14] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][14] ), .ZN(n2330) );
  NAND3_X1 U2357 ( .A1(n2332), .A2(n2331), .A3(n2330), .ZN(n2333) );
  OR3_X1 U2358 ( .A1(n2335), .A2(n2334), .A3(n2333), .ZN(\xmem_inst/N265 ) );
  AOI22_X1 U2359 ( .A1(n3252), .A2(\xmem_inst/mem[15][28] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][28] ), .ZN(n2339) );
  AOI22_X1 U2360 ( .A1(n3573), .A2(\xmem_inst/mem[29][28] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][28] ), .ZN(n2338) );
  AOI22_X1 U2361 ( .A1(n3253), .A2(\xmem_inst/mem[24][28] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][28] ), .ZN(n2337) );
  AOI22_X1 U2362 ( .A1(n3584), .A2(\xmem_inst/mem[20][28] ), .B1(n3628), .B2(
        \xmem_inst/mem[1][28] ), .ZN(n2336) );
  NAND4_X1 U2363 ( .A1(n2339), .A2(n2338), .A3(n2337), .A4(n2336), .ZN(n2355)
         );
  AOI22_X1 U2364 ( .A1(n3597), .A2(\xmem_inst/mem[35][28] ), .B1(n3629), .B2(
        \xmem_inst/mem[31][28] ), .ZN(n2343) );
  AOI22_X1 U2365 ( .A1(n3625), .A2(\xmem_inst/mem[6][28] ), .B1(n3604), .B2(
        \xmem_inst/mem[4][28] ), .ZN(n2342) );
  AOI22_X1 U2366 ( .A1(n3616), .A2(\xmem_inst/mem[14][28] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][28] ), .ZN(n2341) );
  AOI22_X1 U2367 ( .A1(n3594), .A2(\xmem_inst/mem[19][28] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][28] ), .ZN(n2340) );
  NAND4_X1 U2368 ( .A1(n2343), .A2(n2342), .A3(n2341), .A4(n2340), .ZN(n2354)
         );
  AOI22_X1 U2369 ( .A1(n3626), .A2(\xmem_inst/mem[3][28] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][28] ), .ZN(n2347) );
  AOI22_X1 U2370 ( .A1(n3615), .A2(\xmem_inst/mem[2][28] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][28] ), .ZN(n2346) );
  AOI22_X1 U2371 ( .A1(n3233), .A2(\xmem_inst/mem[0][28] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][28] ), .ZN(n2345) );
  AOI22_X1 U2372 ( .A1(n3574), .A2(\xmem_inst/mem[27][28] ), .B1(n3624), .B2(
        \xmem_inst/mem[11][28] ), .ZN(n2344) );
  NAND4_X1 U2373 ( .A1(n2347), .A2(n2346), .A3(n2345), .A4(n2344), .ZN(n2353)
         );
  AOI22_X1 U2374 ( .A1(n3190), .A2(\xmem_inst/mem[41][28] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][28] ), .ZN(n2351) );
  NAND2_X1 U2375 ( .A1(n3245), .A2(\xmem_inst/mem[42][28] ), .ZN(n2350) );
  NAND2_X1 U2376 ( .A1(n3572), .A2(\xmem_inst/mem[25][28] ), .ZN(n2349) );
  NAND2_X1 U2377 ( .A1(n3220), .A2(\xmem_inst/mem[36][28] ), .ZN(n2348) );
  NAND4_X1 U2378 ( .A1(n2351), .A2(n2350), .A3(n2349), .A4(n2348), .ZN(n2352)
         );
  OR4_X1 U2379 ( .A1(n2355), .A2(n2354), .A3(n2353), .A4(n2352), .ZN(n2365) );
  AOI22_X1 U2380 ( .A1(n3627), .A2(\xmem_inst/mem[39][28] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][28] ), .ZN(n2359) );
  AOI22_X1 U2381 ( .A1(n2958), .A2(\xmem_inst/mem[34][28] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][28] ), .ZN(n2358) );
  AOI22_X1 U2382 ( .A1(n3600), .A2(\xmem_inst/mem[21][28] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][28] ), .ZN(n2357) );
  AOI22_X1 U2383 ( .A1(n2967), .A2(\xmem_inst/mem[23][28] ), .B1(n3184), .B2(
        \xmem_inst/mem[37][28] ), .ZN(n2356) );
  NAND4_X1 U2384 ( .A1(n2359), .A2(n2358), .A3(n2357), .A4(n2356), .ZN(n2364)
         );
  AOI22_X1 U2385 ( .A1(n3580), .A2(\xmem_inst/mem[38][28] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][28] ), .ZN(n2362) );
  AOI22_X1 U2386 ( .A1(n3568), .A2(\xmem_inst/mem[18][28] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][28] ), .ZN(n2361) );
  AOI22_X1 U2387 ( .A1(n3148), .A2(\xmem_inst/mem[32][28] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][28] ), .ZN(n2360) );
  NAND3_X1 U2388 ( .A1(n2362), .A2(n2361), .A3(n2360), .ZN(n2363) );
  OR3_X1 U2389 ( .A1(n2365), .A2(n2364), .A3(n2363), .ZN(\xmem_inst/N251 ) );
  AOI22_X1 U2390 ( .A1(n3627), .A2(\xmem_inst/mem[39][9] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][9] ), .ZN(n2369) );
  AOI22_X1 U2391 ( .A1(n3584), .A2(\xmem_inst/mem[20][9] ), .B1(n3602), .B2(
        \xmem_inst/mem[32][9] ), .ZN(n2368) );
  AOI22_X1 U2392 ( .A1(n3580), .A2(\xmem_inst/mem[38][9] ), .B1(n3613), .B2(
        \xmem_inst/mem[37][9] ), .ZN(n2367) );
  AOI22_X1 U2393 ( .A1(n3574), .A2(\xmem_inst/mem[27][9] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][9] ), .ZN(n2366) );
  NAND4_X1 U2394 ( .A1(n2369), .A2(n2368), .A3(n2367), .A4(n2366), .ZN(n2385)
         );
  AOI22_X1 U2395 ( .A1(n3629), .A2(\xmem_inst/mem[31][9] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][9] ), .ZN(n2373) );
  AOI22_X1 U2396 ( .A1(n3624), .A2(\xmem_inst/mem[11][9] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][9] ), .ZN(n2372) );
  AOI22_X1 U2397 ( .A1(n3244), .A2(\xmem_inst/mem[29][9] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][9] ), .ZN(n2371) );
  AOI22_X1 U2398 ( .A1(n3615), .A2(\xmem_inst/mem[2][9] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][9] ), .ZN(n2370) );
  NAND4_X1 U2399 ( .A1(n2373), .A2(n2372), .A3(n2371), .A4(n2370), .ZN(n2384)
         );
  AOI22_X1 U2400 ( .A1(n3235), .A2(\xmem_inst/mem[6][9] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][9] ), .ZN(n2377) );
  AOI22_X1 U2401 ( .A1(n3614), .A2(\xmem_inst/mem[23][9] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][9] ), .ZN(n2376) );
  AOI22_X1 U2402 ( .A1(n3630), .A2(\xmem_inst/mem[30][9] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][9] ), .ZN(n2375) );
  AOI22_X1 U2403 ( .A1(n3233), .A2(\xmem_inst/mem[0][9] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][9] ), .ZN(n2374) );
  NAND4_X1 U2404 ( .A1(n2377), .A2(n2376), .A3(n2375), .A4(n2374), .ZN(n2383)
         );
  AOI22_X1 U2405 ( .A1(n3593), .A2(\xmem_inst/mem[40][9] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][9] ), .ZN(n2381) );
  NAND2_X1 U2406 ( .A1(n3190), .A2(\xmem_inst/mem[41][9] ), .ZN(n2380) );
  NAND2_X1 U2407 ( .A1(n3604), .A2(\xmem_inst/mem[4][9] ), .ZN(n2379) );
  NAND2_X1 U2408 ( .A1(n3220), .A2(\xmem_inst/mem[36][9] ), .ZN(n2378) );
  NAND4_X1 U2409 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n2382)
         );
  OR4_X1 U2410 ( .A1(n2385), .A2(n2384), .A3(n2383), .A4(n2382), .ZN(n2395) );
  AOI22_X1 U2411 ( .A1(n3597), .A2(\xmem_inst/mem[35][9] ), .B1(n3616), .B2(
        \xmem_inst/mem[14][9] ), .ZN(n2389) );
  AOI22_X1 U2412 ( .A1(n3252), .A2(\xmem_inst/mem[15][9] ), .B1(n3572), .B2(
        \xmem_inst/mem[25][9] ), .ZN(n2388) );
  AOI22_X1 U2413 ( .A1(n3628), .A2(\xmem_inst/mem[1][9] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][9] ), .ZN(n2387) );
  AOI22_X1 U2414 ( .A1(n3225), .A2(\xmem_inst/mem[5][9] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][9] ), .ZN(n2386) );
  NAND4_X1 U2415 ( .A1(n2389), .A2(n2388), .A3(n2387), .A4(n2386), .ZN(n2394)
         );
  AOI22_X1 U2416 ( .A1(n3626), .A2(\xmem_inst/mem[3][9] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][9] ), .ZN(n2392) );
  AOI22_X1 U2417 ( .A1(n3568), .A2(\xmem_inst/mem[18][9] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][9] ), .ZN(n2391) );
  AOI22_X1 U2418 ( .A1(n3226), .A2(\xmem_inst/mem[33][9] ), .B1(n3631), .B2(
        \xmem_inst/mem[34][9] ), .ZN(n2390) );
  NAND3_X1 U2419 ( .A1(n2392), .A2(n2391), .A3(n2390), .ZN(n2393) );
  OR3_X1 U2420 ( .A1(n2395), .A2(n2394), .A3(n2393), .ZN(\xmem_inst/N270 ) );
  AOI22_X1 U2421 ( .A1(n3219), .A2(\xmem_inst/mem[9][16] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][16] ), .ZN(n2399) );
  AOI22_X1 U2422 ( .A1(n3613), .A2(\xmem_inst/mem[37][16] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][16] ), .ZN(n2398) );
  AOI22_X1 U2423 ( .A1(n3626), .A2(\xmem_inst/mem[3][16] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][16] ), .ZN(n2397) );
  AOI22_X1 U2424 ( .A1(n3220), .A2(\xmem_inst/mem[36][16] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][16] ), .ZN(n2396) );
  NAND4_X1 U2425 ( .A1(n2399), .A2(n2398), .A3(n2397), .A4(n2396), .ZN(n2415)
         );
  AOI22_X1 U2426 ( .A1(n3233), .A2(\xmem_inst/mem[0][16] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][16] ), .ZN(n2403) );
  AOI22_X1 U2427 ( .A1(n3614), .A2(\xmem_inst/mem[23][16] ), .B1(n3602), .B2(
        \xmem_inst/mem[32][16] ), .ZN(n2402) );
  AOI22_X1 U2428 ( .A1(n3628), .A2(\xmem_inst/mem[1][16] ), .B1(n3572), .B2(
        \xmem_inst/mem[25][16] ), .ZN(n2401) );
  AOI22_X1 U2429 ( .A1(n3604), .A2(\xmem_inst/mem[4][16] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][16] ), .ZN(n2400) );
  NAND4_X1 U2430 ( .A1(n2403), .A2(n2402), .A3(n2401), .A4(n2400), .ZN(n2414)
         );
  AOI22_X1 U2431 ( .A1(n3582), .A2(\xmem_inst/mem[7][16] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][16] ), .ZN(n2407) );
  AOI22_X1 U2432 ( .A1(n3235), .A2(\xmem_inst/mem[6][16] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][16] ), .ZN(n2406) );
  AOI22_X1 U2433 ( .A1(n3580), .A2(\xmem_inst/mem[38][16] ), .B1(n3252), .B2(
        \xmem_inst/mem[15][16] ), .ZN(n2405) );
  AOI22_X1 U2434 ( .A1(n3629), .A2(\xmem_inst/mem[31][16] ), .B1(n3568), .B2(
        \xmem_inst/mem[18][16] ), .ZN(n2404) );
  NAND4_X1 U2435 ( .A1(n2407), .A2(n2406), .A3(n2405), .A4(n2404), .ZN(n2413)
         );
  AOI22_X1 U2436 ( .A1(n3597), .A2(\xmem_inst/mem[35][16] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][16] ), .ZN(n2411) );
  NAND2_X1 U2437 ( .A1(n3617), .A2(\xmem_inst/mem[42][16] ), .ZN(n2410) );
  NAND2_X1 U2438 ( .A1(n3615), .A2(\xmem_inst/mem[2][16] ), .ZN(n2409) );
  NAND2_X1 U2439 ( .A1(n3583), .A2(\xmem_inst/mem[12][16] ), .ZN(n2408) );
  NAND4_X1 U2440 ( .A1(n2411), .A2(n2410), .A3(n2409), .A4(n2408), .ZN(n2412)
         );
  OR4_X1 U2441 ( .A1(n2415), .A2(n2414), .A3(n2413), .A4(n2412), .ZN(n2425) );
  AOI22_X1 U2442 ( .A1(n3586), .A2(\xmem_inst/mem[24][16] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][16] ), .ZN(n2419) );
  AOI22_X1 U2443 ( .A1(n3616), .A2(\xmem_inst/mem[14][16] ), .B1(n3244), .B2(
        \xmem_inst/mem[29][16] ), .ZN(n2418) );
  AOI22_X1 U2444 ( .A1(n3631), .A2(\xmem_inst/mem[34][16] ), .B1(n3574), .B2(
        \xmem_inst/mem[27][16] ), .ZN(n2417) );
  AOI22_X1 U2445 ( .A1(n3627), .A2(\xmem_inst/mem[39][16] ), .B1(n3251), .B2(
        \xmem_inst/mem[20][16] ), .ZN(n2416) );
  NAND4_X1 U2446 ( .A1(n2419), .A2(n2418), .A3(n2417), .A4(n2416), .ZN(n2424)
         );
  AOI22_X1 U2447 ( .A1(n3592), .A2(\xmem_inst/mem[41][16] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][16] ), .ZN(n2422) );
  AOI22_X1 U2448 ( .A1(n3624), .A2(\xmem_inst/mem[11][16] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][16] ), .ZN(n2421) );
  AOI22_X1 U2449 ( .A1(n3569), .A2(\xmem_inst/mem[13][16] ), .B1(n3591), .B2(
        \xmem_inst/mem[8][16] ), .ZN(n2420) );
  NAND3_X1 U2450 ( .A1(n2422), .A2(n2421), .A3(n2420), .ZN(n2423) );
  OR3_X1 U2451 ( .A1(n2425), .A2(n2424), .A3(n2423), .ZN(\xmem_inst/N263 ) );
  AOI22_X1 U2452 ( .A1(n3627), .A2(\xmem_inst/mem[39][13] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][13] ), .ZN(n2429) );
  AOI22_X1 U2453 ( .A1(n3235), .A2(\xmem_inst/mem[6][13] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][13] ), .ZN(n2428) );
  AOI22_X1 U2454 ( .A1(n3584), .A2(\xmem_inst/mem[20][13] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][13] ), .ZN(n2427) );
  AOI22_X1 U2455 ( .A1(n3626), .A2(\xmem_inst/mem[3][13] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][13] ), .ZN(n2426) );
  NAND4_X1 U2456 ( .A1(n2429), .A2(n2428), .A3(n2427), .A4(n2426), .ZN(n2445)
         );
  AOI22_X1 U2457 ( .A1(n3574), .A2(\xmem_inst/mem[27][13] ), .B1(n3604), .B2(
        \xmem_inst/mem[4][13] ), .ZN(n2433) );
  AOI22_X1 U2458 ( .A1(n3233), .A2(\xmem_inst/mem[0][13] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][13] ), .ZN(n2432) );
  AOI22_X1 U2459 ( .A1(n3614), .A2(\xmem_inst/mem[23][13] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][13] ), .ZN(n2431) );
  AOI22_X1 U2460 ( .A1(n3591), .A2(\xmem_inst/mem[8][13] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][13] ), .ZN(n2430) );
  NAND4_X1 U2461 ( .A1(n2433), .A2(n2432), .A3(n2431), .A4(n2430), .ZN(n2444)
         );
  AOI22_X1 U2462 ( .A1(n3244), .A2(\xmem_inst/mem[29][13] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][13] ), .ZN(n2437) );
  NAND2_X1 U2463 ( .A1(n3190), .A2(\xmem_inst/mem[41][13] ), .ZN(n2436) );
  NAND2_X1 U2464 ( .A1(n3582), .A2(\xmem_inst/mem[7][13] ), .ZN(n2435) );
  NAND2_X1 U2465 ( .A1(n3571), .A2(\xmem_inst/mem[28][13] ), .ZN(n2434) );
  AND4_X1 U2466 ( .A1(n2437), .A2(n2436), .A3(n2435), .A4(n2434), .ZN(n2439)
         );
  AOI22_X1 U2467 ( .A1(n3631), .A2(\xmem_inst/mem[34][13] ), .B1(n3580), .B2(
        \xmem_inst/mem[38][13] ), .ZN(n2438) );
  NAND2_X1 U2468 ( .A1(n2439), .A2(n2438), .ZN(n2443) );
  AOI22_X1 U2469 ( .A1(n3629), .A2(\xmem_inst/mem[31][13] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][13] ), .ZN(n2441) );
  AOI22_X1 U2470 ( .A1(n3597), .A2(\xmem_inst/mem[35][13] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][13] ), .ZN(n2440) );
  NAND2_X1 U2471 ( .A1(n2441), .A2(n2440), .ZN(n2442) );
  OR4_X1 U2472 ( .A1(n2445), .A2(n2444), .A3(n2443), .A4(n2442), .ZN(n2456) );
  AOI22_X1 U2473 ( .A1(n3220), .A2(\xmem_inst/mem[36][13] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][13] ), .ZN(n2449) );
  AOI22_X1 U2474 ( .A1(n3586), .A2(\xmem_inst/mem[24][13] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][13] ), .ZN(n2448) );
  AOI22_X1 U2475 ( .A1(n3615), .A2(\xmem_inst/mem[2][13] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][13] ), .ZN(n2447) );
  AOI22_X1 U2476 ( .A1(n3252), .A2(\xmem_inst/mem[15][13] ), .B1(n3184), .B2(
        \xmem_inst/mem[37][13] ), .ZN(n2446) );
  NAND4_X1 U2477 ( .A1(n2449), .A2(n2448), .A3(n2447), .A4(n2446), .ZN(n2455)
         );
  AOI22_X1 U2478 ( .A1(n3568), .A2(\xmem_inst/mem[18][13] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][13] ), .ZN(n2453) );
  AOI22_X1 U2479 ( .A1(n3585), .A2(\xmem_inst/mem[16][13] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][13] ), .ZN(n2452) );
  AOI22_X1 U2480 ( .A1(n3616), .A2(\xmem_inst/mem[14][13] ), .B1(n3624), .B2(
        \xmem_inst/mem[11][13] ), .ZN(n2451) );
  AOI22_X1 U2481 ( .A1(n3602), .A2(\xmem_inst/mem[32][13] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][13] ), .ZN(n2450) );
  NAND4_X1 U2482 ( .A1(n2453), .A2(n2452), .A3(n2451), .A4(n2450), .ZN(n2454)
         );
  OR3_X1 U2483 ( .A1(n2456), .A2(n2455), .A3(n2454), .ZN(\xmem_inst/N266 ) );
  AOI22_X1 U2484 ( .A1(n3628), .A2(\xmem_inst/mem[1][15] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][15] ), .ZN(n2460) );
  AOI22_X1 U2485 ( .A1(n3629), .A2(\xmem_inst/mem[31][15] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][15] ), .ZN(n2459) );
  AOI22_X1 U2486 ( .A1(n3601), .A2(\xmem_inst/mem[26][15] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][15] ), .ZN(n2458) );
  AOI22_X1 U2487 ( .A1(n3616), .A2(\xmem_inst/mem[14][15] ), .B1(n3624), .B2(
        \xmem_inst/mem[11][15] ), .ZN(n2457) );
  NAND4_X1 U2488 ( .A1(n2460), .A2(n2459), .A3(n2458), .A4(n2457), .ZN(n2476)
         );
  AOI22_X1 U2489 ( .A1(n3597), .A2(\xmem_inst/mem[35][15] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][15] ), .ZN(n2464) );
  AOI22_X1 U2490 ( .A1(n3234), .A2(\xmem_inst/mem[2][15] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][15] ), .ZN(n2463) );
  AOI22_X1 U2491 ( .A1(n3613), .A2(\xmem_inst/mem[37][15] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][15] ), .ZN(n2462) );
  AOI22_X1 U2492 ( .A1(n3594), .A2(\xmem_inst/mem[19][15] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][15] ), .ZN(n2461) );
  NAND4_X1 U2493 ( .A1(n2464), .A2(n2463), .A3(n2462), .A4(n2461), .ZN(n2475)
         );
  AOI22_X1 U2494 ( .A1(n3585), .A2(\xmem_inst/mem[16][15] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][15] ), .ZN(n2466) );
  AOI22_X1 U2495 ( .A1(n3574), .A2(\xmem_inst/mem[27][15] ), .B1(n3592), .B2(
        \xmem_inst/mem[41][15] ), .ZN(n2465) );
  NAND2_X1 U2496 ( .A1(n2466), .A2(n2465), .ZN(n2474) );
  AOI22_X1 U2497 ( .A1(\xmem_inst/mem[23][15] ), .A2(n3614), .B1(n3568), .B2(
        \xmem_inst/mem[18][15] ), .ZN(n2470) );
  NAND2_X1 U2498 ( .A1(n2972), .A2(\xmem_inst/mem[40][15] ), .ZN(n2469) );
  NAND2_X1 U2499 ( .A1(n3627), .A2(\xmem_inst/mem[39][15] ), .ZN(n2468) );
  NAND2_X1 U2500 ( .A1(n3631), .A2(\xmem_inst/mem[34][15] ), .ZN(n2467) );
  AND4_X1 U2501 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), .ZN(n2472)
         );
  AOI22_X1 U2502 ( .A1(n3179), .A2(\xmem_inst/mem[8][15] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][15] ), .ZN(n2471) );
  NAND2_X1 U2503 ( .A1(n2472), .A2(n2471), .ZN(n2473) );
  OR4_X1 U2504 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .ZN(n2487) );
  AOI22_X1 U2505 ( .A1(n3096), .A2(\xmem_inst/mem[10][15] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][15] ), .ZN(n2480) );
  AOI22_X1 U2506 ( .A1(n3252), .A2(\xmem_inst/mem[15][15] ), .B1(n3244), .B2(
        \xmem_inst/mem[29][15] ), .ZN(n2479) );
  AOI22_X1 U2507 ( .A1(n3600), .A2(\xmem_inst/mem[21][15] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][15] ), .ZN(n2478) );
  AOI22_X1 U2508 ( .A1(n3625), .A2(\xmem_inst/mem[6][15] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][15] ), .ZN(n2477) );
  NAND4_X1 U2509 ( .A1(n2480), .A2(n2479), .A3(n2478), .A4(n2477), .ZN(n2486)
         );
  AOI22_X1 U2510 ( .A1(n3584), .A2(\xmem_inst/mem[20][15] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][15] ), .ZN(n2484) );
  AOI22_X1 U2511 ( .A1(n3233), .A2(\xmem_inst/mem[0][15] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][15] ), .ZN(n2483) );
  AOI22_X1 U2512 ( .A1(n3586), .A2(\xmem_inst/mem[24][15] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][15] ), .ZN(n2482) );
  AOI22_X1 U2513 ( .A1(n3580), .A2(\xmem_inst/mem[38][15] ), .B1(n3602), .B2(
        \xmem_inst/mem[32][15] ), .ZN(n2481) );
  NAND4_X1 U2514 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n2485)
         );
  OR3_X1 U2515 ( .A1(n2487), .A2(n2486), .A3(n2485), .ZN(\xmem_inst/N264 ) );
  AOI22_X1 U2516 ( .A1(n3573), .A2(\xmem_inst/mem[29][25] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][25] ), .ZN(n2491) );
  AOI22_X1 U2517 ( .A1(n3219), .A2(\xmem_inst/mem[9][25] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][25] ), .ZN(n2490) );
  AOI22_X1 U2518 ( .A1(n3571), .A2(\xmem_inst/mem[28][25] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][25] ), .ZN(n2489) );
  AOI22_X1 U2519 ( .A1(n3624), .A2(\xmem_inst/mem[11][25] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][25] ), .ZN(n2488) );
  NAND4_X1 U2520 ( .A1(n2491), .A2(n2490), .A3(n2489), .A4(n2488), .ZN(n2507)
         );
  AOI22_X1 U2521 ( .A1(n3584), .A2(\xmem_inst/mem[20][25] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][25] ), .ZN(n2495) );
  AOI22_X1 U2522 ( .A1(n3252), .A2(\xmem_inst/mem[15][25] ), .B1(n3572), .B2(
        \xmem_inst/mem[25][25] ), .ZN(n2494) );
  AOI22_X1 U2523 ( .A1(n3580), .A2(\xmem_inst/mem[38][25] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][25] ), .ZN(n2493) );
  AOI22_X1 U2524 ( .A1(n3631), .A2(\xmem_inst/mem[34][25] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][25] ), .ZN(n2492) );
  NAND4_X1 U2525 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n2506)
         );
  AOI22_X1 U2526 ( .A1(n3568), .A2(\xmem_inst/mem[18][25] ), .B1(n3190), .B2(
        \xmem_inst/mem[41][25] ), .ZN(n2497) );
  AOI22_X1 U2527 ( .A1(n3627), .A2(\xmem_inst/mem[39][25] ), .B1(n3617), .B2(
        \xmem_inst/mem[42][25] ), .ZN(n2496) );
  NAND2_X1 U2528 ( .A1(n2497), .A2(n2496), .ZN(n2505) );
  AOI22_X1 U2529 ( .A1(n3616), .A2(\xmem_inst/mem[14][25] ), .B1(n3629), .B2(
        \xmem_inst/mem[31][25] ), .ZN(n2501) );
  NAND2_X1 U2530 ( .A1(n3593), .A2(\xmem_inst/mem[40][25] ), .ZN(n2500) );
  NAND2_X1 U2531 ( .A1(n3582), .A2(\xmem_inst/mem[7][25] ), .ZN(n2499) );
  NAND2_X1 U2532 ( .A1(n3628), .A2(\xmem_inst/mem[1][25] ), .ZN(n2498) );
  AND4_X1 U2533 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n2503)
         );
  AOI22_X1 U2534 ( .A1(n3625), .A2(\xmem_inst/mem[6][25] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][25] ), .ZN(n2502) );
  NAND2_X1 U2535 ( .A1(n2503), .A2(n2502), .ZN(n2504) );
  OR4_X1 U2536 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n2518) );
  AOI22_X1 U2537 ( .A1(n3602), .A2(\xmem_inst/mem[32][25] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][25] ), .ZN(n2511) );
  AOI22_X1 U2538 ( .A1(n3600), .A2(\xmem_inst/mem[21][25] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][25] ), .ZN(n2510) );
  AOI22_X1 U2539 ( .A1(n3084), .A2(\xmem_inst/mem[16][25] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][25] ), .ZN(n2509) );
  AOI22_X1 U2540 ( .A1(n2967), .A2(\xmem_inst/mem[23][25] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][25] ), .ZN(n2508) );
  NAND4_X1 U2541 ( .A1(n2511), .A2(n2510), .A3(n2509), .A4(n2508), .ZN(n2517)
         );
  AOI22_X1 U2542 ( .A1(n3615), .A2(\xmem_inst/mem[2][25] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][25] ), .ZN(n2515) );
  AOI22_X1 U2543 ( .A1(n3233), .A2(\xmem_inst/mem[0][25] ), .B1(n3597), .B2(
        \xmem_inst/mem[35][25] ), .ZN(n2514) );
  AOI22_X1 U2544 ( .A1(n3574), .A2(\xmem_inst/mem[27][25] ), .B1(n3184), .B2(
        \xmem_inst/mem[37][25] ), .ZN(n2513) );
  AOI22_X1 U2545 ( .A1(n3604), .A2(\xmem_inst/mem[4][25] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][25] ), .ZN(n2512) );
  NAND4_X1 U2546 ( .A1(n2515), .A2(n2514), .A3(n2513), .A4(n2512), .ZN(n2516)
         );
  OR3_X1 U2547 ( .A1(n2518), .A2(n2517), .A3(n2516), .ZN(\xmem_inst/N254 ) );
  AOI22_X1 U2548 ( .A1(n3250), .A2(\xmem_inst/mem[27][30] ), .B1(n3613), .B2(
        \xmem_inst/mem[37][30] ), .ZN(n2522) );
  AOI22_X1 U2549 ( .A1(n3628), .A2(\xmem_inst/mem[1][30] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][30] ), .ZN(n2521) );
  AOI22_X1 U2550 ( .A1(n3154), .A2(\xmem_inst/mem[14][30] ), .B1(n3252), .B2(
        \xmem_inst/mem[15][30] ), .ZN(n2520) );
  AOI22_X1 U2551 ( .A1(n3604), .A2(\xmem_inst/mem[4][30] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][30] ), .ZN(n2519) );
  NAND4_X1 U2552 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), .ZN(n2538)
         );
  AOI22_X1 U2553 ( .A1(n3235), .A2(\xmem_inst/mem[6][30] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][30] ), .ZN(n2526) );
  AOI22_X1 U2554 ( .A1(n3220), .A2(\xmem_inst/mem[36][30] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][30] ), .ZN(n2525) );
  AOI22_X1 U2555 ( .A1(n3594), .A2(\xmem_inst/mem[19][30] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][30] ), .ZN(n2524) );
  AOI22_X1 U2556 ( .A1(n3234), .A2(\xmem_inst/mem[2][30] ), .B1(n3580), .B2(
        \xmem_inst/mem[38][30] ), .ZN(n2523) );
  NAND4_X1 U2557 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n2537)
         );
  AOI22_X1 U2558 ( .A1(n3584), .A2(\xmem_inst/mem[20][30] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][30] ), .ZN(n2530) );
  NAND2_X1 U2559 ( .A1(n3190), .A2(\xmem_inst/mem[41][30] ), .ZN(n2529) );
  NAND2_X1 U2560 ( .A1(n3627), .A2(\xmem_inst/mem[39][30] ), .ZN(n2528) );
  NAND2_X1 U2561 ( .A1(n3572), .A2(\xmem_inst/mem[25][30] ), .ZN(n2527) );
  AND4_X1 U2562 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n2532)
         );
  AOI22_X1 U2563 ( .A1(n3614), .A2(\xmem_inst/mem[23][30] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][30] ), .ZN(n2531) );
  NAND2_X1 U2564 ( .A1(n2532), .A2(n2531), .ZN(n2536) );
  AOI22_X1 U2565 ( .A1(n3233), .A2(\xmem_inst/mem[0][30] ), .B1(n3617), .B2(
        \xmem_inst/mem[42][30] ), .ZN(n2534) );
  AOI22_X1 U2566 ( .A1(n3253), .A2(\xmem_inst/mem[24][30] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][30] ), .ZN(n2533) );
  NAND2_X1 U2567 ( .A1(n2534), .A2(n2533), .ZN(n2535) );
  OR4_X1 U2568 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), .ZN(n2549) );
  AOI22_X1 U2569 ( .A1(n3602), .A2(\xmem_inst/mem[32][30] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][30] ), .ZN(n2542) );
  AOI22_X1 U2570 ( .A1(n3626), .A2(\xmem_inst/mem[3][30] ), .B1(n3581), .B2(
        \xmem_inst/mem[22][30] ), .ZN(n2541) );
  AOI22_X1 U2571 ( .A1(n3254), .A2(\xmem_inst/mem[11][30] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][30] ), .ZN(n2540) );
  AOI22_X1 U2572 ( .A1(n3568), .A2(\xmem_inst/mem[18][30] ), .B1(n3573), .B2(
        \xmem_inst/mem[29][30] ), .ZN(n2539) );
  NAND4_X1 U2573 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), .ZN(n2548)
         );
  AOI22_X1 U2574 ( .A1(n2958), .A2(\xmem_inst/mem[34][30] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][30] ), .ZN(n2546) );
  AOI22_X1 U2575 ( .A1(n3597), .A2(\xmem_inst/mem[35][30] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][30] ), .ZN(n2545) );
  AOI22_X1 U2576 ( .A1(n3603), .A2(\xmem_inst/mem[10][30] ), .B1(n3591), .B2(
        \xmem_inst/mem[8][30] ), .ZN(n2544) );
  AOI22_X1 U2577 ( .A1(n3629), .A2(\xmem_inst/mem[31][30] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][30] ), .ZN(n2543) );
  NAND4_X1 U2578 ( .A1(n2546), .A2(n2545), .A3(n2544), .A4(n2543), .ZN(n2547)
         );
  OR3_X1 U2579 ( .A1(n2549), .A2(n2548), .A3(n2547), .ZN(\xmem_inst/N249 ) );
  AOI22_X1 U2580 ( .A1(n3234), .A2(\xmem_inst/mem[2][23] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][23] ), .ZN(n2553) );
  AOI22_X1 U2581 ( .A1(n2967), .A2(\xmem_inst/mem[23][23] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][23] ), .ZN(n2552) );
  AOI22_X1 U2582 ( .A1(n2958), .A2(\xmem_inst/mem[34][23] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][23] ), .ZN(n2551) );
  AOI22_X1 U2583 ( .A1(n3072), .A2(\xmem_inst/mem[31][23] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][23] ), .ZN(n2550) );
  NAND4_X1 U2584 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n2569)
         );
  AOI22_X1 U2585 ( .A1(n3571), .A2(\xmem_inst/mem[28][23] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][23] ), .ZN(n2557) );
  AOI22_X1 U2586 ( .A1(n3233), .A2(\xmem_inst/mem[0][23] ), .B1(n3602), .B2(
        \xmem_inst/mem[32][23] ), .ZN(n2556) );
  AOI22_X1 U2587 ( .A1(n3628), .A2(\xmem_inst/mem[1][23] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][23] ), .ZN(n2555) );
  AOI22_X1 U2588 ( .A1(n3613), .A2(\xmem_inst/mem[37][23] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][23] ), .ZN(n2554) );
  NAND4_X1 U2589 ( .A1(n2557), .A2(n2556), .A3(n2555), .A4(n2554), .ZN(n2568)
         );
  AOI22_X1 U2590 ( .A1(n3580), .A2(\xmem_inst/mem[38][23] ), .B1(n3617), .B2(
        \xmem_inst/mem[42][23] ), .ZN(n2559) );
  AOI22_X1 U2591 ( .A1(n3626), .A2(\xmem_inst/mem[3][23] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][23] ), .ZN(n2558) );
  NAND2_X1 U2592 ( .A1(n2559), .A2(n2558), .ZN(n2567) );
  AOI22_X1 U2593 ( .A1(n3616), .A2(\xmem_inst/mem[14][23] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][23] ), .ZN(n2563) );
  NAND2_X1 U2594 ( .A1(n3190), .A2(\xmem_inst/mem[41][23] ), .ZN(n2562) );
  NAND2_X1 U2595 ( .A1(n3597), .A2(\xmem_inst/mem[35][23] ), .ZN(n2561) );
  NAND2_X1 U2596 ( .A1(n3570), .A2(\xmem_inst/mem[17][23] ), .ZN(n2560) );
  AND4_X1 U2597 ( .A1(n2563), .A2(n2562), .A3(n2561), .A4(n2560), .ZN(n2565)
         );
  AOI22_X1 U2598 ( .A1(n3625), .A2(\xmem_inst/mem[6][23] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][23] ), .ZN(n2564) );
  NAND2_X1 U2599 ( .A1(n2565), .A2(n2564), .ZN(n2566) );
  OR4_X1 U2600 ( .A1(n2569), .A2(n2568), .A3(n2567), .A4(n2566), .ZN(n2580) );
  AOI22_X1 U2601 ( .A1(n3624), .A2(\xmem_inst/mem[11][23] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][23] ), .ZN(n2573) );
  AOI22_X1 U2602 ( .A1(n3153), .A2(\xmem_inst/mem[18][23] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][23] ), .ZN(n2572) );
  AOI22_X1 U2603 ( .A1(n3574), .A2(\xmem_inst/mem[27][23] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][23] ), .ZN(n2571) );
  AOI22_X1 U2604 ( .A1(n3253), .A2(\xmem_inst/mem[24][23] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][23] ), .ZN(n2570) );
  NAND4_X1 U2605 ( .A1(n2573), .A2(n2572), .A3(n2571), .A4(n2570), .ZN(n2579)
         );
  AOI22_X1 U2606 ( .A1(n3584), .A2(\xmem_inst/mem[20][23] ), .B1(n3208), .B2(
        \xmem_inst/mem[26][23] ), .ZN(n2577) );
  AOI22_X1 U2607 ( .A1(n3627), .A2(\xmem_inst/mem[39][23] ), .B1(n3252), .B2(
        \xmem_inst/mem[15][23] ), .ZN(n2576) );
  AOI22_X1 U2608 ( .A1(n3572), .A2(\xmem_inst/mem[25][23] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][23] ), .ZN(n2575) );
  AOI22_X1 U2609 ( .A1(n3244), .A2(\xmem_inst/mem[29][23] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][23] ), .ZN(n2574) );
  NAND4_X1 U2610 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n2578)
         );
  OR3_X1 U2611 ( .A1(n2580), .A2(n2579), .A3(n2578), .ZN(\xmem_inst/N256 ) );
  NOR2_X1 U2612 ( .A1(n4077), .A2(fmem_addr[1]), .ZN(n3690) );
  NOR2_X1 U2613 ( .A1(fmem_addr[0]), .A2(fmem_addr[2]), .ZN(n2582) );
  NOR2_X1 U2614 ( .A1(n3690), .A2(n2582), .ZN(\fmem_inst/N62 ) );
  OR2_X1 U2615 ( .A1(fmem_addr[3]), .A2(fmem_addr[0]), .ZN(n2593) );
  OAI21_X1 U2616 ( .B1(fmem_addr[1]), .B2(fmem_addr[0]), .A(n2593), .ZN(
        \fmem_inst/N75 ) );
  NAND2_X1 U2617 ( .A1(fmem_addr[1]), .A2(fmem_addr[2]), .ZN(n2612) );
  INV_X1 U2618 ( .A(n2612), .ZN(n2590) );
  NAND2_X1 U2619 ( .A1(n2593), .A2(n2590), .ZN(\fmem_inst/N78 ) );
  NAND2_X1 U2620 ( .A1(n4074), .A2(fmem_addr[2]), .ZN(n2594) );
  NOR2_X1 U2621 ( .A1(n3690), .A2(n2594), .ZN(n2589) );
  INV_X1 U2622 ( .A(n2589), .ZN(n2581) );
  AND2_X1 U2623 ( .A1(n4069), .A2(fmem_addr[2]), .ZN(n2606) );
  NAND2_X1 U2624 ( .A1(n2606), .A2(fmem_addr[3]), .ZN(n3695) );
  NAND2_X1 U2625 ( .A1(n4069), .A2(n4078), .ZN(n2600) );
  INV_X1 U2626 ( .A(n2600), .ZN(n2583) );
  AND2_X1 U2627 ( .A1(fmem_addr[3]), .A2(fmem_addr[0]), .ZN(n2585) );
  NAND2_X1 U2628 ( .A1(n2583), .A2(n2585), .ZN(n2592) );
  NAND2_X1 U2629 ( .A1(n4078), .A2(fmem_addr[1]), .ZN(n2595) );
  INV_X1 U2630 ( .A(n2595), .ZN(n2587) );
  NAND2_X1 U2631 ( .A1(n2587), .A2(fmem_addr[3]), .ZN(n3682) );
  NAND4_X1 U2632 ( .A1(n2581), .A2(n3695), .A3(n2592), .A4(n3682), .ZN(
        \fmem_inst/N70 ) );
  NOR2_X1 U2633 ( .A1(n4074), .A2(fmem_addr[3]), .ZN(n3691) );
  NOR3_X1 U2634 ( .A1(n2583), .A2(n3691), .A3(n2582), .ZN(n2584) );
  OAI21_X1 U2635 ( .B1(n4077), .B2(n2612), .A(n2584), .ZN(\fmem_inst/N64 ) );
  NAND2_X1 U2636 ( .A1(n4074), .A2(fmem_addr[3]), .ZN(n2599) );
  NAND2_X1 U2637 ( .A1(n2585), .A2(n2590), .ZN(n4012) );
  NAND2_X1 U2638 ( .A1(n4077), .A2(n4069), .ZN(n2586) );
  OAI211_X1 U2639 ( .C1(fmem_addr[2]), .C2(n2599), .A(n4012), .B(n2586), .ZN(
        \fmem_inst/N69 ) );
  INV_X1 U2640 ( .A(n2593), .ZN(n3689) );
  AOI211_X1 U2641 ( .C1(fmem_addr[1]), .C2(n3689), .A(n3690), .B(n2587), .ZN(
        n2588) );
  NAND2_X1 U2642 ( .A1(n3691), .A2(n2606), .ZN(n3683) );
  NAND2_X1 U2643 ( .A1(n2588), .A2(n3683), .ZN(\fmem_inst/N74 ) );
  OAI22_X1 U2644 ( .A1(n3695), .A2(n4074), .B1(n2595), .B2(n2599), .ZN(n2596)
         );
  NOR2_X1 U2645 ( .A1(n2600), .A2(fmem_addr[0]), .ZN(n3693) );
  NOR3_X1 U2646 ( .A1(n2596), .A2(n3693), .A3(n2589), .ZN(n3686) );
  NAND2_X1 U2647 ( .A1(n3691), .A2(n2590), .ZN(n2591) );
  NAND2_X1 U2648 ( .A1(n3686), .A2(n2591), .ZN(\fmem_inst/N73 ) );
  OAI21_X1 U2649 ( .B1(n2595), .B2(n2593), .A(n2591), .ZN(n2598) );
  INV_X1 U2650 ( .A(n2598), .ZN(n3688) );
  NAND4_X1 U2651 ( .A1(n3688), .A2(n2594), .A3(n2593), .A4(n2592), .ZN(
        \fmem_inst/N63 ) );
  NOR2_X1 U2652 ( .A1(n2595), .A2(n4074), .ZN(n2607) );
  INV_X1 U2653 ( .A(n2607), .ZN(n3685) );
  NAND2_X1 U2654 ( .A1(n3689), .A2(n4069), .ZN(n3684) );
  OAI211_X1 U2655 ( .C1(fmem_addr[3]), .C2(n2600), .A(n3685), .B(n3684), .ZN(
        n2597) );
  OR3_X1 U2656 ( .A1(n2597), .A2(n2596), .A3(n2598), .ZN(\fmem_inst/N72 ) );
  NOR2_X1 U2657 ( .A1(n4097), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[19]) );
  NOR2_X1 U2658 ( .A1(n4098), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[20]) );
  NOR2_X1 U2659 ( .A1(n4095), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[17]) );
  NOR2_X1 U2660 ( .A1(n4096), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[18]) );
  NOR2_X1 U2661 ( .A1(n4101), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[23]) );
  NOR2_X1 U2662 ( .A1(n326), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[24]) );
  NOR2_X1 U2663 ( .A1(n327), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[25]) );
  NOR2_X1 U2664 ( .A1(n328), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[26]) );
  NOR2_X1 U2665 ( .A1(n318), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[27]) );
  NOR2_X1 U2666 ( .A1(n319), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[28]) );
  NOR2_X1 U2667 ( .A1(n4093), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[15]) );
  NOR2_X1 U2668 ( .A1(n4092), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[14]) );
  NOR2_X1 U2669 ( .A1(n4091), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[13]) );
  NOR2_X1 U2670 ( .A1(n4090), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[12]) );
  NOR2_X1 U2671 ( .A1(n325), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[11]) );
  NOR2_X1 U2672 ( .A1(n322), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[10]) );
  NOR2_X1 U2673 ( .A1(n324), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[9]) );
  NOR2_X1 U2674 ( .A1(n323), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[8]) );
  NOR2_X1 U2675 ( .A1(n4089), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[7]) );
  NOR2_X1 U2676 ( .A1(n4088), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[6]) );
  NOR2_X1 U2677 ( .A1(n4104), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[5]) );
  NOR2_X1 U2678 ( .A1(n4103), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[4]) );
  NOR2_X1 U2679 ( .A1(n4087), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[3]) );
  NOR2_X1 U2680 ( .A1(n4086), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[2]) );
  NOR2_X1 U2681 ( .A1(n4085), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[1]) );
  NOR2_X1 U2682 ( .A1(n4084), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[0]) );
  NOR2_X1 U2683 ( .A1(n4099), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[21]) );
  NOR2_X1 U2684 ( .A1(n4100), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[22]) );
  NOR2_X1 U2685 ( .A1(n320), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[29]) );
  NOR2_X1 U2686 ( .A1(n4094), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[16]) );
  NOR2_X1 U2687 ( .A1(n321), .A2(\mac_unit_inst/adder_reg [31]), .ZN(
        m_data_out_y[30]) );
  AOI211_X1 U2688 ( .C1(n2606), .C2(n3689), .A(n2607), .B(n2598), .ZN(n2602)
         );
  OAI21_X1 U2689 ( .B1(n2599), .B2(n2612), .A(n2602), .ZN(\fmem_inst/N65 ) );
  INV_X1 U2690 ( .A(n2606), .ZN(n2603) );
  NOR2_X1 U2691 ( .A1(n2600), .A2(n4077), .ZN(n2601) );
  NOR2_X1 U2692 ( .A1(n2601), .A2(n3691), .ZN(n3687) );
  OAI211_X1 U2693 ( .C1(n4074), .C2(n2603), .A(n2602), .B(n3687), .ZN(
        \fmem_inst/N77 ) );
  NAND3_X1 U2694 ( .A1(n4071), .A2(n4009), .A3(n4010), .ZN(n2619) );
  NOR2_X1 U2695 ( .A1(conv_done), .A2(reset), .ZN(n4025) );
  OAI21_X1 U2696 ( .B1(n2604), .B2(n4009), .A(n4025), .ZN(n2614) );
  NOR2_X1 U2697 ( .A1(n2619), .A2(n4074), .ZN(n2611) );
  OR2_X1 U2698 ( .A1(n2614), .A2(n2611), .ZN(n2610) );
  AOI21_X1 U2699 ( .B1(n2619), .B2(n4074), .A(n2610), .ZN(n104) );
  INV_X1 U2700 ( .A(n2619), .ZN(n2605) );
  OAI21_X1 U2701 ( .B1(n2607), .B2(n2606), .A(n2605), .ZN(n2608) );
  OAI22_X1 U2702 ( .A1(n2610), .A2(n4078), .B1(n2608), .B2(n2614), .ZN(n102)
         );
  NAND2_X1 U2703 ( .A1(n4069), .A2(n2611), .ZN(n2609) );
  OAI22_X1 U2704 ( .A1(n2610), .A2(n4069), .B1(n2614), .B2(n2609), .ZN(n103)
         );
  INV_X1 U2705 ( .A(n2611), .ZN(n2613) );
  NOR2_X1 U2706 ( .A1(n2613), .A2(n2612), .ZN(n2616) );
  INV_X1 U2707 ( .A(n2614), .ZN(n2620) );
  OAI21_X1 U2708 ( .B1(fmem_addr[3]), .B2(n2616), .A(n2620), .ZN(n2615) );
  AOI21_X1 U2709 ( .B1(fmem_addr[3]), .B2(n2616), .A(n2615), .ZN(n105) );
  INV_X1 U2710 ( .A(n4025), .ZN(n2622) );
  NAND4_X1 U2711 ( .A1(xmem_addr[5]), .A2(xmem_addr[1]), .A3(xmem_addr[3]), 
        .A4(n4081), .ZN(n2617) );
  OR3_X1 U2712 ( .A1(xmem_addr[0]), .A2(xmem_addr[2]), .A3(n2617), .ZN(n2618)
         );
  OAI21_X1 U2713 ( .B1(n3697), .B2(n2618), .A(n4025), .ZN(n4026) );
  OAI22_X1 U2714 ( .A1(n2619), .A2(n2622), .B1(n3697), .B2(n4026), .ZN(n4036)
         );
  INV_X1 U2715 ( .A(n4036), .ZN(n4041) );
  NOR2_X1 U2716 ( .A1(xmem_addr[2]), .A2(n4041), .ZN(n2627) );
  NAND2_X1 U2717 ( .A1(xmem_addr[0]), .A2(xmem_addr[1]), .ZN(n4031) );
  INV_X1 U2718 ( .A(n4031), .ZN(n2626) );
  NAND3_X1 U2719 ( .A1(n2620), .A2(n2619), .A3(n3697), .ZN(n4032) );
  OAI221_X1 U2720 ( .B1(n4041), .B2(xmem_addr[1]), .C1(n4041), .C2(
        xmem_addr[0]), .A(n4032), .ZN(n2623) );
  INV_X1 U2721 ( .A(n4009), .ZN(n4006) );
  NAND2_X1 U2722 ( .A1(n4010), .A2(n4006), .ZN(n2621) );
  NOR2_X1 U2723 ( .A1(n2622), .A2(n2621), .ZN(n4042) );
  AOI22_X1 U2724 ( .A1(xmem_addr[2]), .A2(n2623), .B1(n4042), .B2(
        \ctrl_conv_output_inst/cnt_conv [2]), .ZN(n2624) );
  INV_X1 U2725 ( .A(n2624), .ZN(n2625) );
  AOI21_X1 U2726 ( .B1(n2627), .B2(n2626), .A(n2625), .ZN(n4113) );
  AOI22_X1 U2727 ( .A1(n3184), .A2(\xmem_inst/mem[37][24] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][24] ), .ZN(n2631) );
  AOI22_X1 U2728 ( .A1(n2958), .A2(\xmem_inst/mem[34][24] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][24] ), .ZN(n2630) );
  AOI22_X1 U2729 ( .A1(n3233), .A2(\xmem_inst/mem[0][24] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][24] ), .ZN(n2629) );
  AOI22_X1 U2730 ( .A1(n3604), .A2(\xmem_inst/mem[4][24] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][24] ), .ZN(n2628) );
  NAND4_X1 U2731 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n2645)
         );
  AOI22_X1 U2732 ( .A1(n3234), .A2(\xmem_inst/mem[2][24] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][24] ), .ZN(n2635) );
  AOI22_X1 U2733 ( .A1(n3244), .A2(\xmem_inst/mem[29][24] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][24] ), .ZN(n2634) );
  AOI22_X1 U2734 ( .A1(n3569), .A2(\xmem_inst/mem[13][24] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][24] ), .ZN(n2633) );
  AOI22_X1 U2735 ( .A1(n3581), .A2(\xmem_inst/mem[22][24] ), .B1(n3208), .B2(
        \xmem_inst/mem[26][24] ), .ZN(n2632) );
  NAND4_X1 U2736 ( .A1(n2635), .A2(n2634), .A3(n2633), .A4(n2632), .ZN(n2644)
         );
  AOI22_X1 U2737 ( .A1(n2967), .A2(\xmem_inst/mem[23][24] ), .B1(n3072), .B2(
        \xmem_inst/mem[31][24] ), .ZN(n2639) );
  AOI22_X1 U2738 ( .A1(n3627), .A2(\xmem_inst/mem[39][24] ), .B1(n3624), .B2(
        \xmem_inst/mem[11][24] ), .ZN(n2638) );
  AOI22_X1 U2739 ( .A1(n3572), .A2(\xmem_inst/mem[25][24] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][24] ), .ZN(n2637) );
  AOI22_X1 U2740 ( .A1(n3580), .A2(\xmem_inst/mem[38][24] ), .B1(n3252), .B2(
        \xmem_inst/mem[15][24] ), .ZN(n2636) );
  NAND4_X1 U2741 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .ZN(n2643)
         );
  AOI22_X1 U2742 ( .A1(n3592), .A2(\xmem_inst/mem[41][24] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][24] ), .ZN(n2641) );
  AOI22_X1 U2743 ( .A1(n3153), .A2(\xmem_inst/mem[18][24] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][24] ), .ZN(n2640) );
  NAND2_X1 U2744 ( .A1(n2641), .A2(n2640), .ZN(n2642) );
  NOR4_X1 U2745 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .ZN(n2657)
         );
  AOI22_X1 U2746 ( .A1(n3597), .A2(\xmem_inst/mem[35][24] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][24] ), .ZN(n2656) );
  AOI22_X1 U2747 ( .A1(n3586), .A2(\xmem_inst/mem[24][24] ), .B1(n3616), .B2(
        \xmem_inst/mem[14][24] ), .ZN(n2649) );
  NAND2_X1 U2748 ( .A1(n3593), .A2(\xmem_inst/mem[40][24] ), .ZN(n2648) );
  NAND2_X1 U2749 ( .A1(n3574), .A2(\xmem_inst/mem[27][24] ), .ZN(n2647) );
  NAND2_X1 U2750 ( .A1(n3225), .A2(\xmem_inst/mem[5][24] ), .ZN(n2646) );
  AND4_X1 U2751 ( .A1(n2649), .A2(n2648), .A3(n2647), .A4(n2646), .ZN(n2655)
         );
  AOI22_X1 U2752 ( .A1(n3584), .A2(\xmem_inst/mem[20][24] ), .B1(n3220), .B2(
        \xmem_inst/mem[36][24] ), .ZN(n2653) );
  AOI22_X1 U2753 ( .A1(n3619), .A2(\xmem_inst/mem[9][24] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][24] ), .ZN(n2652) );
  AOI22_X1 U2754 ( .A1(n3602), .A2(\xmem_inst/mem[32][24] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][24] ), .ZN(n2651) );
  AOI22_X1 U2755 ( .A1(n3625), .A2(\xmem_inst/mem[6][24] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][24] ), .ZN(n2650) );
  AND4_X1 U2756 ( .A1(n2653), .A2(n2652), .A3(n2651), .A4(n2650), .ZN(n2654)
         );
  NAND4_X1 U2757 ( .A1(n2657), .A2(n2656), .A3(n2655), .A4(n2654), .ZN(
        \xmem_inst/N255 ) );
  AOI22_X1 U2758 ( .A1(n3627), .A2(\xmem_inst/mem[39][10] ), .B1(n3603), .B2(
        \xmem_inst/mem[10][10] ), .ZN(n2661) );
  AOI22_X1 U2759 ( .A1(n3594), .A2(\xmem_inst/mem[19][10] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][10] ), .ZN(n2660) );
  AOI22_X1 U2760 ( .A1(n3250), .A2(\xmem_inst/mem[27][10] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][10] ), .ZN(n2659) );
  AOI22_X1 U2761 ( .A1(n3254), .A2(\xmem_inst/mem[11][10] ), .B1(n3219), .B2(
        \xmem_inst/mem[9][10] ), .ZN(n2658) );
  NAND4_X1 U2762 ( .A1(n2661), .A2(n2660), .A3(n2659), .A4(n2658), .ZN(n2675)
         );
  AOI22_X1 U2763 ( .A1(n3584), .A2(\xmem_inst/mem[20][10] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][10] ), .ZN(n2665) );
  AOI22_X1 U2764 ( .A1(n3614), .A2(\xmem_inst/mem[23][10] ), .B1(n3220), .B2(
        \xmem_inst/mem[36][10] ), .ZN(n2664) );
  AOI22_X1 U2765 ( .A1(n3598), .A2(\xmem_inst/mem[0][10] ), .B1(n3252), .B2(
        \xmem_inst/mem[15][10] ), .ZN(n2663) );
  AOI22_X1 U2766 ( .A1(n3625), .A2(\xmem_inst/mem[6][10] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][10] ), .ZN(n2662) );
  NAND4_X1 U2767 ( .A1(n2665), .A2(n2664), .A3(n2663), .A4(n2662), .ZN(n2674)
         );
  AOI22_X1 U2768 ( .A1(n3630), .A2(\xmem_inst/mem[30][10] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][10] ), .ZN(n2669) );
  AOI22_X1 U2769 ( .A1(n3615), .A2(\xmem_inst/mem[2][10] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][10] ), .ZN(n2668) );
  AOI22_X1 U2770 ( .A1(n3203), .A2(\xmem_inst/mem[38][10] ), .B1(n3072), .B2(
        \xmem_inst/mem[31][10] ), .ZN(n2667) );
  AOI22_X1 U2771 ( .A1(n3084), .A2(\xmem_inst/mem[16][10] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][10] ), .ZN(n2666) );
  NAND4_X1 U2772 ( .A1(n2669), .A2(n2668), .A3(n2667), .A4(n2666), .ZN(n2673)
         );
  AOI22_X1 U2773 ( .A1(n3613), .A2(\xmem_inst/mem[37][10] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][10] ), .ZN(n2671) );
  AOI22_X1 U2774 ( .A1(n3631), .A2(\xmem_inst/mem[34][10] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][10] ), .ZN(n2670) );
  NAND2_X1 U2775 ( .A1(n2671), .A2(n2670), .ZN(n2672) );
  NOR4_X1 U2776 ( .A1(n2675), .A2(n2674), .A3(n2673), .A4(n2672), .ZN(n2687)
         );
  AOI22_X1 U2777 ( .A1(n3626), .A2(\xmem_inst/mem[3][10] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][10] ), .ZN(n2686) );
  AOI22_X1 U2778 ( .A1(n3244), .A2(\xmem_inst/mem[29][10] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][10] ), .ZN(n2679) );
  NAND2_X1 U2779 ( .A1(n3190), .A2(\xmem_inst/mem[41][10] ), .ZN(n2678) );
  NAND2_X1 U2780 ( .A1(n3597), .A2(\xmem_inst/mem[35][10] ), .ZN(n2677) );
  NAND2_X1 U2781 ( .A1(n3602), .A2(\xmem_inst/mem[32][10] ), .ZN(n2676) );
  AND4_X1 U2782 ( .A1(n2679), .A2(n2678), .A3(n2677), .A4(n2676), .ZN(n2685)
         );
  AOI22_X1 U2783 ( .A1(n3570), .A2(\xmem_inst/mem[17][10] ), .B1(n3599), .B2(
        \xmem_inst/mem[33][10] ), .ZN(n2683) );
  AOI22_X1 U2784 ( .A1(n3628), .A2(\xmem_inst/mem[1][10] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][10] ), .ZN(n2682) );
  AOI22_X1 U2785 ( .A1(n3568), .A2(\xmem_inst/mem[18][10] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][10] ), .ZN(n2681) );
  AOI22_X1 U2786 ( .A1(n3616), .A2(\xmem_inst/mem[14][10] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][10] ), .ZN(n2680) );
  AND4_X1 U2787 ( .A1(n2683), .A2(n2682), .A3(n2681), .A4(n2680), .ZN(n2684)
         );
  NAND4_X1 U2788 ( .A1(n2687), .A2(n2686), .A3(n2685), .A4(n2684), .ZN(
        \xmem_inst/N269 ) );
  AOI22_X1 U2789 ( .A1(n3631), .A2(\xmem_inst/mem[34][2] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][2] ), .ZN(n2691) );
  AOI22_X1 U2790 ( .A1(n3597), .A2(\xmem_inst/mem[35][2] ), .B1(n3599), .B2(
        \xmem_inst/mem[33][2] ), .ZN(n2690) );
  AOI22_X1 U2791 ( .A1(n3604), .A2(\xmem_inst/mem[4][2] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][2] ), .ZN(n2689) );
  AOI22_X1 U2792 ( .A1(n3628), .A2(\xmem_inst/mem[1][2] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][2] ), .ZN(n2688) );
  NAND4_X1 U2793 ( .A1(n2691), .A2(n2690), .A3(n2689), .A4(n2688), .ZN(n2705)
         );
  AOI22_X1 U2794 ( .A1(n3629), .A2(\xmem_inst/mem[31][2] ), .B1(n3153), .B2(
        \xmem_inst/mem[18][2] ), .ZN(n2695) );
  AOI22_X1 U2795 ( .A1(n3614), .A2(\xmem_inst/mem[23][2] ), .B1(n3184), .B2(
        \xmem_inst/mem[37][2] ), .ZN(n2694) );
  AOI22_X1 U2796 ( .A1(n3252), .A2(\xmem_inst/mem[15][2] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][2] ), .ZN(n2693) );
  AOI22_X1 U2797 ( .A1(n3591), .A2(\xmem_inst/mem[8][2] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][2] ), .ZN(n2692) );
  NAND4_X1 U2798 ( .A1(n2695), .A2(n2694), .A3(n2693), .A4(n2692), .ZN(n2704)
         );
  AOI22_X1 U2799 ( .A1(n3253), .A2(\xmem_inst/mem[24][2] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][2] ), .ZN(n2699) );
  AOI22_X1 U2800 ( .A1(n3250), .A2(\xmem_inst/mem[27][2] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][2] ), .ZN(n2698) );
  AOI22_X1 U2801 ( .A1(n3585), .A2(\xmem_inst/mem[16][2] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][2] ), .ZN(n2697) );
  AOI22_X1 U2802 ( .A1(n3235), .A2(\xmem_inst/mem[6][2] ), .B1(n3616), .B2(
        \xmem_inst/mem[14][2] ), .ZN(n2696) );
  NAND4_X1 U2803 ( .A1(n2699), .A2(n2698), .A3(n2697), .A4(n2696), .ZN(n2703)
         );
  AOI22_X1 U2804 ( .A1(n3225), .A2(\xmem_inst/mem[5][2] ), .B1(n3581), .B2(
        \xmem_inst/mem[22][2] ), .ZN(n2701) );
  AOI22_X1 U2805 ( .A1(n3244), .A2(\xmem_inst/mem[29][2] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][2] ), .ZN(n2700) );
  NAND2_X1 U2806 ( .A1(n2701), .A2(n2700), .ZN(n2702) );
  NOR4_X1 U2807 ( .A1(n2705), .A2(n2704), .A3(n2703), .A4(n2702), .ZN(n2717)
         );
  AOI22_X1 U2808 ( .A1(n3593), .A2(\xmem_inst/mem[40][2] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][2] ), .ZN(n2716) );
  AOI22_X1 U2809 ( .A1(n3584), .A2(\xmem_inst/mem[20][2] ), .B1(n3233), .B2(
        \xmem_inst/mem[0][2] ), .ZN(n2709) );
  NAND2_X1 U2810 ( .A1(n3190), .A2(\xmem_inst/mem[41][2] ), .ZN(n2708) );
  NAND2_X1 U2811 ( .A1(n3096), .A2(\xmem_inst/mem[10][2] ), .ZN(n2707) );
  NAND2_X1 U2812 ( .A1(n3602), .A2(\xmem_inst/mem[32][2] ), .ZN(n2706) );
  AND4_X1 U2813 ( .A1(n2709), .A2(n2708), .A3(n2707), .A4(n2706), .ZN(n2715)
         );
  AOI22_X1 U2814 ( .A1(n3627), .A2(\xmem_inst/mem[39][2] ), .B1(n3624), .B2(
        \xmem_inst/mem[11][2] ), .ZN(n2713) );
  AOI22_X1 U2815 ( .A1(n3615), .A2(\xmem_inst/mem[2][2] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][2] ), .ZN(n2712) );
  AOI22_X1 U2816 ( .A1(n3619), .A2(\xmem_inst/mem[9][2] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][2] ), .ZN(n2711) );
  AOI22_X1 U2817 ( .A1(n3203), .A2(\xmem_inst/mem[38][2] ), .B1(n3572), .B2(
        \xmem_inst/mem[25][2] ), .ZN(n2710) );
  AND4_X1 U2818 ( .A1(n2713), .A2(n2712), .A3(n2711), .A4(n2710), .ZN(n2714)
         );
  NAND4_X1 U2819 ( .A1(n2717), .A2(n2716), .A3(n2715), .A4(n2714), .ZN(
        \xmem_inst/N277 ) );
  AOI22_X1 U2820 ( .A1(n3625), .A2(\xmem_inst/mem[6][19] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][19] ), .ZN(n2721) );
  AOI22_X1 U2821 ( .A1(n3602), .A2(\xmem_inst/mem[32][19] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][19] ), .ZN(n2720) );
  AOI22_X1 U2822 ( .A1(n3233), .A2(\xmem_inst/mem[0][19] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][19] ), .ZN(n2719) );
  AOI22_X1 U2823 ( .A1(n2967), .A2(\xmem_inst/mem[23][19] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][19] ), .ZN(n2718) );
  NAND4_X1 U2824 ( .A1(n2721), .A2(n2720), .A3(n2719), .A4(n2718), .ZN(n2735)
         );
  AOI22_X1 U2825 ( .A1(n3244), .A2(\xmem_inst/mem[29][19] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][19] ), .ZN(n2725) );
  AOI22_X1 U2826 ( .A1(n3597), .A2(\xmem_inst/mem[35][19] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][19] ), .ZN(n2724) );
  AOI22_X1 U2827 ( .A1(n3624), .A2(\xmem_inst/mem[11][19] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][19] ), .ZN(n2723) );
  AOI22_X1 U2828 ( .A1(n3154), .A2(\xmem_inst/mem[14][19] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][19] ), .ZN(n2722) );
  NAND4_X1 U2829 ( .A1(n2725), .A2(n2724), .A3(n2723), .A4(n2722), .ZN(n2734)
         );
  AOI22_X1 U2830 ( .A1(n3580), .A2(\xmem_inst/mem[38][19] ), .B1(n3072), .B2(
        \xmem_inst/mem[31][19] ), .ZN(n2729) );
  AOI22_X1 U2831 ( .A1(n3584), .A2(\xmem_inst/mem[20][19] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][19] ), .ZN(n2728) );
  AOI22_X1 U2832 ( .A1(n3604), .A2(\xmem_inst/mem[4][19] ), .B1(n3208), .B2(
        \xmem_inst/mem[26][19] ), .ZN(n2727) );
  AOI22_X1 U2833 ( .A1(n3220), .A2(\xmem_inst/mem[36][19] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][19] ), .ZN(n2726) );
  NAND4_X1 U2834 ( .A1(n2729), .A2(n2728), .A3(n2727), .A4(n2726), .ZN(n2733)
         );
  AOI22_X1 U2835 ( .A1(n3253), .A2(\xmem_inst/mem[24][19] ), .B1(n3190), .B2(
        \xmem_inst/mem[41][19] ), .ZN(n2731) );
  AOI22_X1 U2836 ( .A1(n3568), .A2(\xmem_inst/mem[18][19] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][19] ), .ZN(n2730) );
  NAND2_X1 U2837 ( .A1(n2731), .A2(n2730), .ZN(n2732) );
  NOR4_X1 U2838 ( .A1(n2735), .A2(n2734), .A3(n2733), .A4(n2732), .ZN(n2747)
         );
  AOI22_X1 U2839 ( .A1(n3569), .A2(\xmem_inst/mem[13][19] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][19] ), .ZN(n2746) );
  AOI22_X1 U2840 ( .A1(n3572), .A2(\xmem_inst/mem[25][19] ), .B1(n3250), .B2(
        \xmem_inst/mem[27][19] ), .ZN(n2739) );
  NAND2_X1 U2841 ( .A1(n3593), .A2(\xmem_inst/mem[40][19] ), .ZN(n2738) );
  NAND2_X1 U2842 ( .A1(n3618), .A2(\xmem_inst/mem[15][19] ), .ZN(n2737) );
  NAND2_X1 U2843 ( .A1(n3613), .A2(\xmem_inst/mem[37][19] ), .ZN(n2736) );
  AND4_X1 U2844 ( .A1(n2739), .A2(n2738), .A3(n2737), .A4(n2736), .ZN(n2745)
         );
  AOI22_X1 U2845 ( .A1(n2958), .A2(\xmem_inst/mem[34][19] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][19] ), .ZN(n2743) );
  AOI22_X1 U2846 ( .A1(n3627), .A2(\xmem_inst/mem[39][19] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][19] ), .ZN(n2742) );
  AOI22_X1 U2847 ( .A1(n3615), .A2(\xmem_inst/mem[2][19] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][19] ), .ZN(n2741) );
  AOI22_X1 U2848 ( .A1(n3582), .A2(\xmem_inst/mem[7][19] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][19] ), .ZN(n2740) );
  AND4_X1 U2849 ( .A1(n2743), .A2(n2742), .A3(n2741), .A4(n2740), .ZN(n2744)
         );
  NAND4_X1 U2850 ( .A1(n2747), .A2(n2746), .A3(n2745), .A4(n2744), .ZN(
        \xmem_inst/N260 ) );
  AOI22_X1 U2851 ( .A1(n3631), .A2(\xmem_inst/mem[34][3] ), .B1(n3251), .B2(
        \xmem_inst/mem[20][3] ), .ZN(n2751) );
  AOI22_X1 U2852 ( .A1(n3203), .A2(\xmem_inst/mem[38][3] ), .B1(n3624), .B2(
        \xmem_inst/mem[11][3] ), .ZN(n2750) );
  AOI22_X1 U2853 ( .A1(n3625), .A2(\xmem_inst/mem[6][3] ), .B1(n3153), .B2(
        \xmem_inst/mem[18][3] ), .ZN(n2749) );
  AOI22_X1 U2854 ( .A1(n3084), .A2(\xmem_inst/mem[16][3] ), .B1(n3219), .B2(
        \xmem_inst/mem[9][3] ), .ZN(n2748) );
  NAND4_X1 U2855 ( .A1(n2751), .A2(n2750), .A3(n2749), .A4(n2748), .ZN(n2765)
         );
  AOI22_X1 U2856 ( .A1(n3627), .A2(\xmem_inst/mem[39][3] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][3] ), .ZN(n2755) );
  AOI22_X1 U2857 ( .A1(n3629), .A2(\xmem_inst/mem[31][3] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][3] ), .ZN(n2754) );
  AOI22_X1 U2858 ( .A1(n3148), .A2(\xmem_inst/mem[32][3] ), .B1(n3581), .B2(
        \xmem_inst/mem[22][3] ), .ZN(n2753) );
  AOI22_X1 U2859 ( .A1(n3613), .A2(\xmem_inst/mem[37][3] ), .B1(n3572), .B2(
        \xmem_inst/mem[25][3] ), .ZN(n2752) );
  NAND4_X1 U2860 ( .A1(n2755), .A2(n2754), .A3(n2753), .A4(n2752), .ZN(n2764)
         );
  AOI22_X1 U2861 ( .A1(n3600), .A2(\xmem_inst/mem[21][3] ), .B1(n3604), .B2(
        \xmem_inst/mem[4][3] ), .ZN(n2759) );
  AOI22_X1 U2862 ( .A1(n3225), .A2(\xmem_inst/mem[5][3] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][3] ), .ZN(n2758) );
  AOI22_X1 U2863 ( .A1(n3250), .A2(\xmem_inst/mem[27][3] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][3] ), .ZN(n2757) );
  AOI22_X1 U2864 ( .A1(n3614), .A2(\xmem_inst/mem[23][3] ), .B1(n3597), .B2(
        \xmem_inst/mem[35][3] ), .ZN(n2756) );
  NAND4_X1 U2865 ( .A1(n2759), .A2(n2758), .A3(n2757), .A4(n2756), .ZN(n2763)
         );
  AOI22_X1 U2866 ( .A1(n3598), .A2(\xmem_inst/mem[0][3] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][3] ), .ZN(n2761) );
  AOI22_X1 U2867 ( .A1(n3616), .A2(\xmem_inst/mem[14][3] ), .B1(n3190), .B2(
        \xmem_inst/mem[41][3] ), .ZN(n2760) );
  NAND2_X1 U2868 ( .A1(n2761), .A2(n2760), .ZN(n2762) );
  NOR4_X1 U2869 ( .A1(n2765), .A2(n2764), .A3(n2763), .A4(n2762), .ZN(n2777)
         );
  AOI22_X1 U2870 ( .A1(n3593), .A2(\xmem_inst/mem[40][3] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][3] ), .ZN(n2776) );
  AOI22_X1 U2871 ( .A1(n3571), .A2(\xmem_inst/mem[28][3] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][3] ), .ZN(n2769) );
  NAND2_X1 U2872 ( .A1(n3617), .A2(\xmem_inst/mem[42][3] ), .ZN(n2768) );
  NAND2_X1 U2873 ( .A1(n3626), .A2(\xmem_inst/mem[3][3] ), .ZN(n2767) );
  NAND2_X1 U2874 ( .A1(n3226), .A2(\xmem_inst/mem[33][3] ), .ZN(n2766) );
  AND4_X1 U2875 ( .A1(n2769), .A2(n2768), .A3(n2767), .A4(n2766), .ZN(n2775)
         );
  AOI22_X1 U2876 ( .A1(n3615), .A2(\xmem_inst/mem[2][3] ), .B1(n3220), .B2(
        \xmem_inst/mem[36][3] ), .ZN(n2773) );
  AOI22_X1 U2877 ( .A1(n3244), .A2(\xmem_inst/mem[29][3] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][3] ), .ZN(n2772) );
  AOI22_X1 U2878 ( .A1(n3252), .A2(\xmem_inst/mem[15][3] ), .B1(n3628), .B2(
        \xmem_inst/mem[1][3] ), .ZN(n2771) );
  AOI22_X1 U2879 ( .A1(n3594), .A2(\xmem_inst/mem[19][3] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][3] ), .ZN(n2770) );
  AND4_X1 U2880 ( .A1(n2773), .A2(n2772), .A3(n2771), .A4(n2770), .ZN(n2774)
         );
  NAND4_X1 U2881 ( .A1(n2777), .A2(n2776), .A3(n2775), .A4(n2774), .ZN(
        \xmem_inst/N276 ) );
  AOI22_X1 U2882 ( .A1(n3618), .A2(\xmem_inst/mem[15][26] ), .B1(n3184), .B2(
        \xmem_inst/mem[37][26] ), .ZN(n2781) );
  AOI22_X1 U2883 ( .A1(n3626), .A2(\xmem_inst/mem[3][26] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][26] ), .ZN(n2780) );
  AOI22_X1 U2884 ( .A1(n3574), .A2(\xmem_inst/mem[27][26] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][26] ), .ZN(n2779) );
  AOI22_X1 U2885 ( .A1(n3625), .A2(\xmem_inst/mem[6][26] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][26] ), .ZN(n2778) );
  NAND4_X1 U2886 ( .A1(n2781), .A2(n2780), .A3(n2779), .A4(n2778), .ZN(n2795)
         );
  AOI22_X1 U2887 ( .A1(n3627), .A2(\xmem_inst/mem[39][26] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][26] ), .ZN(n2785) );
  AOI22_X1 U2888 ( .A1(n3154), .A2(\xmem_inst/mem[14][26] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][26] ), .ZN(n2784) );
  AOI22_X1 U2889 ( .A1(n3569), .A2(\xmem_inst/mem[13][26] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][26] ), .ZN(n2783) );
  AOI22_X1 U2890 ( .A1(n3603), .A2(\xmem_inst/mem[10][26] ), .B1(n3208), .B2(
        \xmem_inst/mem[26][26] ), .ZN(n2782) );
  NAND4_X1 U2891 ( .A1(n2785), .A2(n2784), .A3(n2783), .A4(n2782), .ZN(n2794)
         );
  AOI22_X1 U2892 ( .A1(n3580), .A2(\xmem_inst/mem[38][26] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][26] ), .ZN(n2789) );
  AOI22_X1 U2893 ( .A1(n3072), .A2(\xmem_inst/mem[31][26] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][26] ), .ZN(n2788) );
  AOI22_X1 U2894 ( .A1(n3584), .A2(\xmem_inst/mem[20][26] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][26] ), .ZN(n2787) );
  AOI22_X1 U2895 ( .A1(n3234), .A2(\xmem_inst/mem[2][26] ), .B1(n3573), .B2(
        \xmem_inst/mem[29][26] ), .ZN(n2786) );
  NAND4_X1 U2896 ( .A1(n2789), .A2(n2788), .A3(n2787), .A4(n2786), .ZN(n2793)
         );
  AOI22_X1 U2897 ( .A1(n2958), .A2(\xmem_inst/mem[34][26] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][26] ), .ZN(n2791) );
  AOI22_X1 U2898 ( .A1(n3233), .A2(\xmem_inst/mem[0][26] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][26] ), .ZN(n2790) );
  NAND2_X1 U2899 ( .A1(n2791), .A2(n2790), .ZN(n2792) );
  NOR4_X1 U2900 ( .A1(n2795), .A2(n2794), .A3(n2793), .A4(n2792), .ZN(n2807)
         );
  AOI22_X1 U2901 ( .A1(n3592), .A2(\xmem_inst/mem[41][26] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][26] ), .ZN(n2806) );
  AOI22_X1 U2902 ( .A1(n3179), .A2(\xmem_inst/mem[8][26] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][26] ), .ZN(n2799) );
  NAND2_X1 U2903 ( .A1(n3593), .A2(\xmem_inst/mem[40][26] ), .ZN(n2798) );
  NAND2_X1 U2904 ( .A1(n3624), .A2(\xmem_inst/mem[11][26] ), .ZN(n2797) );
  NAND2_X1 U2905 ( .A1(n3225), .A2(\xmem_inst/mem[5][26] ), .ZN(n2796) );
  AND4_X1 U2906 ( .A1(n2799), .A2(n2798), .A3(n2797), .A4(n2796), .ZN(n2805)
         );
  AOI22_X1 U2907 ( .A1(n2967), .A2(\xmem_inst/mem[23][26] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][26] ), .ZN(n2803) );
  AOI22_X1 U2908 ( .A1(n3597), .A2(\xmem_inst/mem[35][26] ), .B1(n3153), .B2(
        \xmem_inst/mem[18][26] ), .ZN(n2802) );
  AOI22_X1 U2909 ( .A1(n3602), .A2(\xmem_inst/mem[32][26] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][26] ), .ZN(n2801) );
  AOI22_X1 U2910 ( .A1(n3600), .A2(\xmem_inst/mem[21][26] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][26] ), .ZN(n2800) );
  AND4_X1 U2911 ( .A1(n2803), .A2(n2802), .A3(n2801), .A4(n2800), .ZN(n2804)
         );
  NAND4_X1 U2912 ( .A1(n2807), .A2(n2806), .A3(n2805), .A4(n2804), .ZN(
        \xmem_inst/N253 ) );
  AOI22_X1 U2913 ( .A1(n3220), .A2(\xmem_inst/mem[36][22] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][22] ), .ZN(n2811) );
  AOI22_X1 U2914 ( .A1(n3625), .A2(\xmem_inst/mem[6][22] ), .B1(n3234), .B2(
        \xmem_inst/mem[2][22] ), .ZN(n2810) );
  AOI22_X1 U2915 ( .A1(n3627), .A2(\xmem_inst/mem[39][22] ), .B1(n3184), .B2(
        \xmem_inst/mem[37][22] ), .ZN(n2809) );
  AOI22_X1 U2916 ( .A1(n3624), .A2(\xmem_inst/mem[11][22] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][22] ), .ZN(n2808) );
  NAND4_X1 U2917 ( .A1(n2811), .A2(n2810), .A3(n2809), .A4(n2808), .ZN(n2825)
         );
  AOI22_X1 U2918 ( .A1(n3601), .A2(\xmem_inst/mem[26][22] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][22] ), .ZN(n2815) );
  AOI22_X1 U2919 ( .A1(n3244), .A2(\xmem_inst/mem[29][22] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][22] ), .ZN(n2814) );
  AOI22_X1 U2920 ( .A1(n3574), .A2(\xmem_inst/mem[27][22] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][22] ), .ZN(n2813) );
  AOI22_X1 U2921 ( .A1(n3580), .A2(\xmem_inst/mem[38][22] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][22] ), .ZN(n2812) );
  NAND4_X1 U2922 ( .A1(n2815), .A2(n2814), .A3(n2813), .A4(n2812), .ZN(n2824)
         );
  AOI22_X1 U2923 ( .A1(n3591), .A2(\xmem_inst/mem[8][22] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][22] ), .ZN(n2819) );
  AOI22_X1 U2924 ( .A1(n3594), .A2(\xmem_inst/mem[19][22] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][22] ), .ZN(n2818) );
  AOI22_X1 U2925 ( .A1(n3154), .A2(\xmem_inst/mem[14][22] ), .B1(n3604), .B2(
        \xmem_inst/mem[4][22] ), .ZN(n2817) );
  AOI22_X1 U2926 ( .A1(n2958), .A2(\xmem_inst/mem[34][22] ), .B1(n3614), .B2(
        \xmem_inst/mem[23][22] ), .ZN(n2816) );
  NAND4_X1 U2927 ( .A1(n2819), .A2(n2818), .A3(n2817), .A4(n2816), .ZN(n2823)
         );
  AOI22_X1 U2928 ( .A1(n3253), .A2(\xmem_inst/mem[24][22] ), .B1(n3190), .B2(
        \xmem_inst/mem[41][22] ), .ZN(n2821) );
  AOI22_X1 U2929 ( .A1(n3597), .A2(\xmem_inst/mem[35][22] ), .B1(n3593), .B2(
        \xmem_inst/mem[40][22] ), .ZN(n2820) );
  NAND2_X1 U2930 ( .A1(n2821), .A2(n2820), .ZN(n2822) );
  NOR4_X1 U2931 ( .A1(n2825), .A2(n2824), .A3(n2823), .A4(n2822), .ZN(n2837)
         );
  AOI22_X1 U2932 ( .A1(n3629), .A2(\xmem_inst/mem[31][22] ), .B1(n3602), .B2(
        \xmem_inst/mem[32][22] ), .ZN(n2836) );
  AOI22_X1 U2933 ( .A1(n3584), .A2(\xmem_inst/mem[20][22] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][22] ), .ZN(n2829) );
  NAND2_X1 U2934 ( .A1(n3245), .A2(\xmem_inst/mem[42][22] ), .ZN(n2828) );
  NAND2_X1 U2935 ( .A1(n3618), .A2(\xmem_inst/mem[15][22] ), .ZN(n2827) );
  NAND2_X1 U2936 ( .A1(n3585), .A2(\xmem_inst/mem[16][22] ), .ZN(n2826) );
  AND4_X1 U2937 ( .A1(n2829), .A2(n2828), .A3(n2827), .A4(n2826), .ZN(n2835)
         );
  AOI22_X1 U2938 ( .A1(n3600), .A2(\xmem_inst/mem[21][22] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][22] ), .ZN(n2833) );
  AOI22_X1 U2939 ( .A1(n3568), .A2(\xmem_inst/mem[18][22] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][22] ), .ZN(n2832) );
  AOI22_X1 U2940 ( .A1(n3233), .A2(\xmem_inst/mem[0][22] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][22] ), .ZN(n2831) );
  AOI22_X1 U2941 ( .A1(n3096), .A2(\xmem_inst/mem[10][22] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][22] ), .ZN(n2830) );
  AND4_X1 U2942 ( .A1(n2833), .A2(n2832), .A3(n2831), .A4(n2830), .ZN(n2834)
         );
  NAND4_X1 U2943 ( .A1(n2837), .A2(n2836), .A3(n2835), .A4(n2834), .ZN(
        \xmem_inst/N257 ) );
  AOI22_X1 U2944 ( .A1(n3618), .A2(\xmem_inst/mem[15][29] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][29] ), .ZN(n2841) );
  AOI22_X1 U2945 ( .A1(n3233), .A2(\xmem_inst/mem[0][29] ), .B1(n3153), .B2(
        \xmem_inst/mem[18][29] ), .ZN(n2840) );
  AOI22_X1 U2946 ( .A1(n3597), .A2(\xmem_inst/mem[35][29] ), .B1(n3604), .B2(
        \xmem_inst/mem[4][29] ), .ZN(n2839) );
  AOI22_X1 U2947 ( .A1(n3570), .A2(\xmem_inst/mem[17][29] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][29] ), .ZN(n2838) );
  NAND4_X1 U2948 ( .A1(n2841), .A2(n2840), .A3(n2839), .A4(n2838), .ZN(n2855)
         );
  AOI22_X1 U2949 ( .A1(n3574), .A2(\xmem_inst/mem[27][29] ), .B1(n3602), .B2(
        \xmem_inst/mem[32][29] ), .ZN(n2845) );
  AOI22_X1 U2950 ( .A1(n3626), .A2(\xmem_inst/mem[3][29] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][29] ), .ZN(n2844) );
  AOI22_X1 U2951 ( .A1(n2958), .A2(\xmem_inst/mem[34][29] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][29] ), .ZN(n2843) );
  AOI22_X1 U2952 ( .A1(n3072), .A2(\xmem_inst/mem[31][29] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][29] ), .ZN(n2842) );
  NAND4_X1 U2953 ( .A1(n2845), .A2(n2844), .A3(n2843), .A4(n2842), .ZN(n2854)
         );
  AOI22_X1 U2954 ( .A1(n3184), .A2(\xmem_inst/mem[37][29] ), .B1(n3603), .B2(
        \xmem_inst/mem[10][29] ), .ZN(n2849) );
  AOI22_X1 U2955 ( .A1(n3225), .A2(\xmem_inst/mem[5][29] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][29] ), .ZN(n2848) );
  AOI22_X1 U2956 ( .A1(n3220), .A2(\xmem_inst/mem[36][29] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][29] ), .ZN(n2847) );
  AOI22_X1 U2957 ( .A1(n3251), .A2(\xmem_inst/mem[20][29] ), .B1(n3573), .B2(
        \xmem_inst/mem[29][29] ), .ZN(n2846) );
  NAND4_X1 U2958 ( .A1(n2849), .A2(n2848), .A3(n2847), .A4(n2846), .ZN(n2853)
         );
  AOI22_X1 U2959 ( .A1(n3592), .A2(\xmem_inst/mem[41][29] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][29] ), .ZN(n2851) );
  AOI22_X1 U2960 ( .A1(n3245), .A2(\xmem_inst/mem[42][29] ), .B1(n3208), .B2(
        \xmem_inst/mem[26][29] ), .ZN(n2850) );
  NAND2_X1 U2961 ( .A1(n2851), .A2(n2850), .ZN(n2852) );
  NOR4_X1 U2962 ( .A1(n2855), .A2(n2854), .A3(n2853), .A4(n2852), .ZN(n2867)
         );
  AOI22_X1 U2963 ( .A1(n3616), .A2(\xmem_inst/mem[14][29] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][29] ), .ZN(n2866) );
  AOI22_X1 U2964 ( .A1(n3586), .A2(\xmem_inst/mem[24][29] ), .B1(n3615), .B2(
        \xmem_inst/mem[2][29] ), .ZN(n2859) );
  NAND2_X1 U2965 ( .A1(n3593), .A2(\xmem_inst/mem[40][29] ), .ZN(n2858) );
  NAND2_X1 U2966 ( .A1(n3254), .A2(\xmem_inst/mem[11][29] ), .ZN(n2857) );
  NAND2_X1 U2967 ( .A1(n3572), .A2(\xmem_inst/mem[25][29] ), .ZN(n2856) );
  AND4_X1 U2968 ( .A1(n2859), .A2(n2858), .A3(n2857), .A4(n2856), .ZN(n2865)
         );
  AOI22_X1 U2969 ( .A1(n3627), .A2(\xmem_inst/mem[39][29] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][29] ), .ZN(n2863) );
  AOI22_X1 U2970 ( .A1(n2967), .A2(\xmem_inst/mem[23][29] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][29] ), .ZN(n2862) );
  AOI22_X1 U2971 ( .A1(n3580), .A2(\xmem_inst/mem[38][29] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][29] ), .ZN(n2861) );
  AOI22_X1 U2972 ( .A1(n3625), .A2(\xmem_inst/mem[6][29] ), .B1(n3628), .B2(
        \xmem_inst/mem[1][29] ), .ZN(n2860) );
  AND4_X1 U2973 ( .A1(n2863), .A2(n2862), .A3(n2861), .A4(n2860), .ZN(n2864)
         );
  NAND4_X1 U2974 ( .A1(n2867), .A2(n2866), .A3(n2865), .A4(n2864), .ZN(
        \xmem_inst/N250 ) );
  AOI22_X1 U2975 ( .A1(n3601), .A2(\xmem_inst/mem[26][27] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][27] ), .ZN(n2871) );
  AOI22_X1 U2976 ( .A1(n3618), .A2(\xmem_inst/mem[15][27] ), .B1(n3602), .B2(
        \xmem_inst/mem[32][27] ), .ZN(n2870) );
  AOI22_X1 U2977 ( .A1(n3234), .A2(\xmem_inst/mem[2][27] ), .B1(n3580), .B2(
        \xmem_inst/mem[38][27] ), .ZN(n2869) );
  AOI22_X1 U2978 ( .A1(n3084), .A2(\xmem_inst/mem[16][27] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][27] ), .ZN(n2868) );
  NAND4_X1 U2979 ( .A1(n2871), .A2(n2870), .A3(n2869), .A4(n2868), .ZN(n2887)
         );
  AOI22_X1 U2980 ( .A1(n3594), .A2(\xmem_inst/mem[19][27] ), .B1(n3220), .B2(
        \xmem_inst/mem[36][27] ), .ZN(n2875) );
  AOI22_X1 U2981 ( .A1(n3625), .A2(\xmem_inst/mem[6][27] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][27] ), .ZN(n2874) );
  AOI22_X1 U2982 ( .A1(n3251), .A2(\xmem_inst/mem[20][27] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][27] ), .ZN(n2873) );
  AOI22_X1 U2983 ( .A1(n3154), .A2(\xmem_inst/mem[14][27] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][27] ), .ZN(n2872) );
  NAND4_X1 U2984 ( .A1(n2875), .A2(n2874), .A3(n2873), .A4(n2872), .ZN(n2886)
         );
  AOI22_X1 U2985 ( .A1(n3573), .A2(\xmem_inst/mem[29][27] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][27] ), .ZN(n2879) );
  AOI22_X1 U2986 ( .A1(n3597), .A2(\xmem_inst/mem[35][27] ), .B1(n3153), .B2(
        \xmem_inst/mem[18][27] ), .ZN(n2878) );
  AOI22_X1 U2987 ( .A1(n3571), .A2(\xmem_inst/mem[28][27] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][27] ), .ZN(n2877) );
  AOI22_X1 U2988 ( .A1(n2967), .A2(\xmem_inst/mem[23][27] ), .B1(n3572), .B2(
        \xmem_inst/mem[25][27] ), .ZN(n2876) );
  NAND4_X1 U2989 ( .A1(n2879), .A2(n2878), .A3(n2877), .A4(n2876), .ZN(n2885)
         );
  AOI22_X1 U2990 ( .A1(n3627), .A2(\xmem_inst/mem[39][27] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][27] ), .ZN(n2883) );
  AOI22_X1 U2991 ( .A1(n3600), .A2(\xmem_inst/mem[21][27] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][27] ), .ZN(n2882) );
  AOI22_X1 U2992 ( .A1(n3574), .A2(\xmem_inst/mem[27][27] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][27] ), .ZN(n2881) );
  AOI22_X1 U2993 ( .A1(n3233), .A2(\xmem_inst/mem[0][27] ), .B1(n3629), .B2(
        \xmem_inst/mem[31][27] ), .ZN(n2880) );
  NAND4_X1 U2994 ( .A1(n2883), .A2(n2882), .A3(n2881), .A4(n2880), .ZN(n2884)
         );
  NOR4_X1 U2995 ( .A1(n2887), .A2(n2886), .A3(n2885), .A4(n2884), .ZN(n2897)
         );
  AOI22_X1 U2996 ( .A1(n3631), .A2(\xmem_inst/mem[34][27] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][27] ), .ZN(n2896) );
  AOI22_X1 U2997 ( .A1(n3583), .A2(\xmem_inst/mem[12][27] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][27] ), .ZN(n2891) );
  NAND2_X1 U2998 ( .A1(n3190), .A2(\xmem_inst/mem[41][27] ), .ZN(n2890) );
  NAND2_X1 U2999 ( .A1(n3254), .A2(\xmem_inst/mem[11][27] ), .ZN(n2889) );
  NAND2_X1 U3000 ( .A1(n3613), .A2(\xmem_inst/mem[37][27] ), .ZN(n2888) );
  AND4_X1 U3001 ( .A1(n2891), .A2(n2890), .A3(n2889), .A4(n2888), .ZN(n2895)
         );
  AOI22_X1 U3002 ( .A1(n3617), .A2(\xmem_inst/mem[42][27] ), .B1(n3628), .B2(
        \xmem_inst/mem[1][27] ), .ZN(n2893) );
  AOI22_X1 U3003 ( .A1(n3570), .A2(\xmem_inst/mem[17][27] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][27] ), .ZN(n2892) );
  AND2_X1 U3004 ( .A1(n2893), .A2(n2892), .ZN(n2894) );
  NAND4_X1 U3005 ( .A1(n2897), .A2(n2896), .A3(n2895), .A4(n2894), .ZN(
        \xmem_inst/N252 ) );
  AOI22_X1 U3006 ( .A1(n3628), .A2(\xmem_inst/mem[1][11] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][11] ), .ZN(n2901) );
  AOI22_X1 U3007 ( .A1(n3148), .A2(\xmem_inst/mem[32][11] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][11] ), .ZN(n2900) );
  AOI22_X1 U3008 ( .A1(n3625), .A2(\xmem_inst/mem[6][11] ), .B1(n3251), .B2(
        \xmem_inst/mem[20][11] ), .ZN(n2899) );
  AOI22_X1 U3009 ( .A1(n3586), .A2(\xmem_inst/mem[24][11] ), .B1(n3581), .B2(
        \xmem_inst/mem[22][11] ), .ZN(n2898) );
  NAND4_X1 U3010 ( .A1(n2901), .A2(n2900), .A3(n2899), .A4(n2898), .ZN(n2915)
         );
  AOI22_X1 U3011 ( .A1(n3203), .A2(\xmem_inst/mem[38][11] ), .B1(n3154), .B2(
        \xmem_inst/mem[14][11] ), .ZN(n2903) );
  AOI22_X1 U3012 ( .A1(n3593), .A2(\xmem_inst/mem[40][11] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][11] ), .ZN(n2902) );
  NAND2_X1 U3013 ( .A1(n2903), .A2(n2902), .ZN(n2914) );
  AOI22_X1 U3014 ( .A1(n3629), .A2(\xmem_inst/mem[31][11] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][11] ), .ZN(n2907) );
  AOI22_X1 U3015 ( .A1(n3613), .A2(\xmem_inst/mem[37][11] ), .B1(n3219), .B2(
        \xmem_inst/mem[9][11] ), .ZN(n2906) );
  AOI22_X1 U3016 ( .A1(n3585), .A2(\xmem_inst/mem[16][11] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][11] ), .ZN(n2905) );
  AOI22_X1 U3017 ( .A1(n3254), .A2(\xmem_inst/mem[11][11] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][11] ), .ZN(n2904) );
  NAND4_X1 U3018 ( .A1(n2907), .A2(n2906), .A3(n2905), .A4(n2904), .ZN(n2913)
         );
  AOI22_X1 U3019 ( .A1(n3252), .A2(\xmem_inst/mem[15][11] ), .B1(n3568), .B2(
        \xmem_inst/mem[18][11] ), .ZN(n2911) );
  AOI22_X1 U3020 ( .A1(n3598), .A2(\xmem_inst/mem[0][11] ), .B1(n3597), .B2(
        \xmem_inst/mem[35][11] ), .ZN(n2910) );
  AOI22_X1 U3021 ( .A1(n3614), .A2(\xmem_inst/mem[23][11] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][11] ), .ZN(n2909) );
  AOI22_X1 U3022 ( .A1(n3631), .A2(\xmem_inst/mem[34][11] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][11] ), .ZN(n2908) );
  NAND4_X1 U3023 ( .A1(n2911), .A2(n2910), .A3(n2909), .A4(n2908), .ZN(n2912)
         );
  NOR4_X1 U3024 ( .A1(n2915), .A2(n2914), .A3(n2913), .A4(n2912), .ZN(n2927)
         );
  AOI22_X1 U3025 ( .A1(n3617), .A2(\xmem_inst/mem[42][11] ), .B1(n3572), .B2(
        \xmem_inst/mem[25][11] ), .ZN(n2926) );
  AOI22_X1 U3026 ( .A1(n3583), .A2(\xmem_inst/mem[12][11] ), .B1(n3250), .B2(
        \xmem_inst/mem[27][11] ), .ZN(n2919) );
  NAND2_X1 U3027 ( .A1(n3190), .A2(\xmem_inst/mem[41][11] ), .ZN(n2918) );
  NAND2_X1 U3028 ( .A1(n3627), .A2(\xmem_inst/mem[39][11] ), .ZN(n2917) );
  NAND2_X1 U3029 ( .A1(n3179), .A2(\xmem_inst/mem[8][11] ), .ZN(n2916) );
  AND4_X1 U3030 ( .A1(n2919), .A2(n2918), .A3(n2917), .A4(n2916), .ZN(n2925)
         );
  AOI22_X1 U3031 ( .A1(n3604), .A2(\xmem_inst/mem[4][11] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][11] ), .ZN(n2923) );
  AOI22_X1 U3032 ( .A1(n3615), .A2(\xmem_inst/mem[2][11] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][11] ), .ZN(n2922) );
  AOI22_X1 U3033 ( .A1(n3244), .A2(\xmem_inst/mem[29][11] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][11] ), .ZN(n2921) );
  AOI22_X1 U3034 ( .A1(n3225), .A2(\xmem_inst/mem[5][11] ), .B1(n3599), .B2(
        \xmem_inst/mem[33][11] ), .ZN(n2920) );
  AND4_X1 U3035 ( .A1(n2923), .A2(n2922), .A3(n2921), .A4(n2920), .ZN(n2924)
         );
  NAND4_X1 U3036 ( .A1(n2927), .A2(n2926), .A3(n2925), .A4(n2924), .ZN(
        \xmem_inst/N268 ) );
  AOI22_X1 U3037 ( .A1(n3072), .A2(\xmem_inst/mem[31][18] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][18] ), .ZN(n2931) );
  AOI22_X1 U3038 ( .A1(n2958), .A2(\xmem_inst/mem[34][18] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][18] ), .ZN(n2930) );
  AOI22_X1 U3039 ( .A1(n3627), .A2(\xmem_inst/mem[39][18] ), .B1(n3208), .B2(
        \xmem_inst/mem[26][18] ), .ZN(n2929) );
  AOI22_X1 U3040 ( .A1(n3618), .A2(\xmem_inst/mem[15][18] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][18] ), .ZN(n2928) );
  NAND4_X1 U3041 ( .A1(n2931), .A2(n2930), .A3(n2929), .A4(n2928), .ZN(n2945)
         );
  AOI22_X1 U3042 ( .A1(n3084), .A2(\xmem_inst/mem[16][18] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][18] ), .ZN(n2935) );
  AOI22_X1 U3043 ( .A1(n3614), .A2(\xmem_inst/mem[23][18] ), .B1(n3251), .B2(
        \xmem_inst/mem[20][18] ), .ZN(n2934) );
  AOI22_X1 U3044 ( .A1(n3154), .A2(\xmem_inst/mem[14][18] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][18] ), .ZN(n2933) );
  AOI22_X1 U3045 ( .A1(n3572), .A2(\xmem_inst/mem[25][18] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][18] ), .ZN(n2932) );
  NAND4_X1 U3046 ( .A1(n2935), .A2(n2934), .A3(n2933), .A4(n2932), .ZN(n2944)
         );
  AOI22_X1 U3047 ( .A1(n3602), .A2(\xmem_inst/mem[32][18] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][18] ), .ZN(n2939) );
  AOI22_X1 U3048 ( .A1(n3597), .A2(\xmem_inst/mem[35][18] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][18] ), .ZN(n2938) );
  AOI22_X1 U3049 ( .A1(n3600), .A2(\xmem_inst/mem[21][18] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][18] ), .ZN(n2937) );
  AOI22_X1 U3050 ( .A1(n3624), .A2(\xmem_inst/mem[11][18] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][18] ), .ZN(n2936) );
  NAND4_X1 U3051 ( .A1(n2939), .A2(n2938), .A3(n2937), .A4(n2936), .ZN(n2943)
         );
  AOI22_X1 U3052 ( .A1(n3244), .A2(\xmem_inst/mem[29][18] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][18] ), .ZN(n2941) );
  AOI22_X1 U3053 ( .A1(n3235), .A2(\xmem_inst/mem[6][18] ), .B1(n3190), .B2(
        \xmem_inst/mem[41][18] ), .ZN(n2940) );
  NAND2_X1 U3054 ( .A1(n2941), .A2(n2940), .ZN(n2942) );
  NOR4_X1 U3055 ( .A1(n2945), .A2(n2944), .A3(n2943), .A4(n2942), .ZN(n2957)
         );
  AOI22_X1 U3056 ( .A1(n3582), .A2(\xmem_inst/mem[7][18] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][18] ), .ZN(n2956) );
  AOI22_X1 U3057 ( .A1(n3253), .A2(\xmem_inst/mem[24][18] ), .B1(n3203), .B2(
        \xmem_inst/mem[38][18] ), .ZN(n2949) );
  NAND2_X1 U3058 ( .A1(n3245), .A2(\xmem_inst/mem[42][18] ), .ZN(n2948) );
  NAND2_X1 U3059 ( .A1(n3615), .A2(\xmem_inst/mem[2][18] ), .ZN(n2947) );
  NAND2_X1 U3060 ( .A1(n3613), .A2(\xmem_inst/mem[37][18] ), .ZN(n2946) );
  AND4_X1 U3061 ( .A1(n2949), .A2(n2948), .A3(n2947), .A4(n2946), .ZN(n2955)
         );
  AOI22_X1 U3062 ( .A1(n3233), .A2(\xmem_inst/mem[0][18] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][18] ), .ZN(n2953) );
  AOI22_X1 U3063 ( .A1(n3568), .A2(\xmem_inst/mem[18][18] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][18] ), .ZN(n2952) );
  AOI22_X1 U3064 ( .A1(n3574), .A2(\xmem_inst/mem[27][18] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][18] ), .ZN(n2951) );
  AOI22_X1 U3065 ( .A1(n3220), .A2(\xmem_inst/mem[36][18] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][18] ), .ZN(n2950) );
  AND4_X1 U3066 ( .A1(n2953), .A2(n2952), .A3(n2951), .A4(n2950), .ZN(n2954)
         );
  NAND4_X1 U3067 ( .A1(n2957), .A2(n2956), .A3(n2955), .A4(n2954), .ZN(
        \xmem_inst/N261 ) );
  AOI22_X1 U3068 ( .A1(n3574), .A2(\xmem_inst/mem[27][21] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][21] ), .ZN(n2962) );
  AOI22_X1 U3069 ( .A1(n3597), .A2(\xmem_inst/mem[35][21] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][21] ), .ZN(n2961) );
  AOI22_X1 U3070 ( .A1(n3219), .A2(\xmem_inst/mem[9][21] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][21] ), .ZN(n2960) );
  AOI22_X1 U3071 ( .A1(n2958), .A2(\xmem_inst/mem[34][21] ), .B1(n3252), .B2(
        \xmem_inst/mem[15][21] ), .ZN(n2959) );
  NAND4_X1 U3072 ( .A1(n2962), .A2(n2961), .A3(n2960), .A4(n2959), .ZN(n2978)
         );
  AOI22_X1 U3073 ( .A1(n3253), .A2(\xmem_inst/mem[24][21] ), .B1(n3153), .B2(
        \xmem_inst/mem[18][21] ), .ZN(n2966) );
  AOI22_X1 U3074 ( .A1(n3154), .A2(\xmem_inst/mem[14][21] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][21] ), .ZN(n2965) );
  AOI22_X1 U3075 ( .A1(n3580), .A2(\xmem_inst/mem[38][21] ), .B1(n3251), .B2(
        \xmem_inst/mem[20][21] ), .ZN(n2964) );
  AOI22_X1 U3076 ( .A1(n3630), .A2(\xmem_inst/mem[30][21] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][21] ), .ZN(n2963) );
  NAND4_X1 U3077 ( .A1(n2966), .A2(n2965), .A3(n2964), .A4(n2963), .ZN(n2977)
         );
  AOI22_X1 U3078 ( .A1(n2967), .A2(\xmem_inst/mem[23][21] ), .B1(n3220), .B2(
        \xmem_inst/mem[36][21] ), .ZN(n2971) );
  AOI22_X1 U3079 ( .A1(n3234), .A2(\xmem_inst/mem[2][21] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][21] ), .ZN(n2970) );
  AOI22_X1 U3080 ( .A1(n3591), .A2(\xmem_inst/mem[8][21] ), .B1(n3208), .B2(
        \xmem_inst/mem[26][21] ), .ZN(n2969) );
  AOI22_X1 U3081 ( .A1(n3625), .A2(\xmem_inst/mem[6][21] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][21] ), .ZN(n2968) );
  NAND4_X1 U3082 ( .A1(n2971), .A2(n2970), .A3(n2969), .A4(n2968), .ZN(n2976)
         );
  AOI22_X1 U3083 ( .A1(n3592), .A2(\xmem_inst/mem[41][21] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][21] ), .ZN(n2974) );
  AOI22_X1 U3084 ( .A1(n3600), .A2(\xmem_inst/mem[21][21] ), .B1(n2972), .B2(
        \xmem_inst/mem[40][21] ), .ZN(n2973) );
  NAND2_X1 U3085 ( .A1(n2974), .A2(n2973), .ZN(n2975) );
  NOR4_X1 U3086 ( .A1(n2978), .A2(n2977), .A3(n2976), .A4(n2975), .ZN(n2990)
         );
  AOI22_X1 U3087 ( .A1(n3613), .A2(\xmem_inst/mem[37][21] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][21] ), .ZN(n2989) );
  AOI22_X1 U3088 ( .A1(n3244), .A2(\xmem_inst/mem[29][21] ), .B1(n3233), .B2(
        \xmem_inst/mem[0][21] ), .ZN(n2982) );
  NAND2_X1 U3089 ( .A1(n3245), .A2(\xmem_inst/mem[42][21] ), .ZN(n2981) );
  NAND2_X1 U3090 ( .A1(n3624), .A2(\xmem_inst/mem[11][21] ), .ZN(n2980) );
  NAND2_X1 U3091 ( .A1(n3225), .A2(\xmem_inst/mem[5][21] ), .ZN(n2979) );
  AND4_X1 U3092 ( .A1(n2982), .A2(n2981), .A3(n2980), .A4(n2979), .ZN(n2988)
         );
  AOI22_X1 U3093 ( .A1(n3594), .A2(\xmem_inst/mem[19][21] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][21] ), .ZN(n2986) );
  AOI22_X1 U3094 ( .A1(n3602), .A2(\xmem_inst/mem[32][21] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][21] ), .ZN(n2985) );
  AOI22_X1 U3095 ( .A1(n3627), .A2(\xmem_inst/mem[39][21] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][21] ), .ZN(n2984) );
  AOI22_X1 U3096 ( .A1(n3072), .A2(\xmem_inst/mem[31][21] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][21] ), .ZN(n2983) );
  AND4_X1 U3097 ( .A1(n2986), .A2(n2985), .A3(n2984), .A4(n2983), .ZN(n2987)
         );
  NAND4_X1 U3098 ( .A1(n2990), .A2(n2989), .A3(n2988), .A4(n2987), .ZN(
        \xmem_inst/N258 ) );
  AOI22_X1 U3099 ( .A1(n3613), .A2(\xmem_inst/mem[37][17] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][17] ), .ZN(n2994) );
  AOI22_X1 U3100 ( .A1(n3084), .A2(\xmem_inst/mem[16][17] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][17] ), .ZN(n2993) );
  AOI22_X1 U3101 ( .A1(n3233), .A2(\xmem_inst/mem[0][17] ), .B1(n3573), .B2(
        \xmem_inst/mem[29][17] ), .ZN(n2992) );
  AOI22_X1 U3102 ( .A1(n3616), .A2(\xmem_inst/mem[14][17] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][17] ), .ZN(n2991) );
  NAND4_X1 U3103 ( .A1(n2994), .A2(n2993), .A3(n2992), .A4(n2991), .ZN(n3010)
         );
  AOI22_X1 U3104 ( .A1(n3597), .A2(\xmem_inst/mem[35][17] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][17] ), .ZN(n2998) );
  AOI22_X1 U3105 ( .A1(n3618), .A2(\xmem_inst/mem[15][17] ), .B1(n3208), .B2(
        \xmem_inst/mem[26][17] ), .ZN(n2997) );
  AOI22_X1 U3106 ( .A1(n3624), .A2(\xmem_inst/mem[11][17] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][17] ), .ZN(n2996) );
  AOI22_X1 U3107 ( .A1(n3572), .A2(\xmem_inst/mem[25][17] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][17] ), .ZN(n2995) );
  NAND4_X1 U3108 ( .A1(n2998), .A2(n2997), .A3(n2996), .A4(n2995), .ZN(n3009)
         );
  AOI22_X1 U3109 ( .A1(n3234), .A2(\xmem_inst/mem[2][17] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][17] ), .ZN(n3002) );
  AOI22_X1 U3110 ( .A1(n3594), .A2(\xmem_inst/mem[19][17] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][17] ), .ZN(n3001) );
  AOI22_X1 U3111 ( .A1(n3627), .A2(\xmem_inst/mem[39][17] ), .B1(n3629), .B2(
        \xmem_inst/mem[31][17] ), .ZN(n3000) );
  AOI22_X1 U3112 ( .A1(n3568), .A2(\xmem_inst/mem[18][17] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][17] ), .ZN(n2999) );
  NAND4_X1 U3113 ( .A1(n3002), .A2(n3001), .A3(n3000), .A4(n2999), .ZN(n3008)
         );
  AOI22_X1 U3114 ( .A1(n3584), .A2(\xmem_inst/mem[20][17] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][17] ), .ZN(n3006) );
  AOI22_X1 U3115 ( .A1(n3604), .A2(\xmem_inst/mem[4][17] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][17] ), .ZN(n3005) );
  AOI22_X1 U3116 ( .A1(n3574), .A2(\xmem_inst/mem[27][17] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][17] ), .ZN(n3004) );
  AOI22_X1 U3117 ( .A1(n3614), .A2(\xmem_inst/mem[23][17] ), .B1(n3625), .B2(
        \xmem_inst/mem[6][17] ), .ZN(n3003) );
  NAND4_X1 U3118 ( .A1(n3006), .A2(n3005), .A3(n3004), .A4(n3003), .ZN(n3007)
         );
  NOR4_X1 U3119 ( .A1(n3010), .A2(n3009), .A3(n3008), .A4(n3007), .ZN(n3019)
         );
  AOI22_X1 U3120 ( .A1(n3617), .A2(\xmem_inst/mem[42][17] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][17] ), .ZN(n3018) );
  AOI22_X1 U3121 ( .A1(n3631), .A2(\xmem_inst/mem[34][17] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][17] ), .ZN(n3017) );
  AOI22_X1 U3122 ( .A1(n3593), .A2(\xmem_inst/mem[40][17] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][17] ), .ZN(n3015) );
  AOI22_X1 U3123 ( .A1(n3602), .A2(\xmem_inst/mem[32][17] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][17] ), .ZN(n3014) );
  AND2_X1 U3124 ( .A1(n3190), .A2(\xmem_inst/mem[41][17] ), .ZN(n3011) );
  AOI21_X1 U3125 ( .B1(n3580), .B2(\xmem_inst/mem[38][17] ), .A(n3011), .ZN(
        n3013) );
  NAND2_X1 U3126 ( .A1(n3220), .A2(\xmem_inst/mem[36][17] ), .ZN(n3012) );
  AND4_X1 U3127 ( .A1(n3015), .A2(n3014), .A3(n3013), .A4(n3012), .ZN(n3016)
         );
  NAND4_X1 U3128 ( .A1(n3019), .A2(n3018), .A3(n3017), .A4(n3016), .ZN(
        \xmem_inst/N262 ) );
  NAND2_X1 U3129 ( .A1(n3617), .A2(\xmem_inst/mem[42][12] ), .ZN(n3020) );
  OAI21_X1 U3130 ( .B1(n3021), .B2(n4107), .A(n3020), .ZN(n3022) );
  AOI21_X1 U3131 ( .B1(n3148), .B2(\xmem_inst/mem[32][12] ), .A(n3022), .ZN(
        n3025) );
  AOI22_X1 U3132 ( .A1(n3614), .A2(\xmem_inst/mem[23][12] ), .B1(n3593), .B2(
        \xmem_inst/mem[40][12] ), .ZN(n3024) );
  AOI22_X1 U3133 ( .A1(n3244), .A2(\xmem_inst/mem[29][12] ), .B1(n3581), .B2(
        \xmem_inst/mem[22][12] ), .ZN(n3023) );
  NAND3_X1 U3134 ( .A1(n3025), .A2(n3024), .A3(n3023), .ZN(n3041) );
  AOI22_X1 U3135 ( .A1(n3604), .A2(\xmem_inst/mem[4][12] ), .B1(n3599), .B2(
        \xmem_inst/mem[33][12] ), .ZN(n3029) );
  AOI22_X1 U3136 ( .A1(n3219), .A2(\xmem_inst/mem[9][12] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][12] ), .ZN(n3028) );
  AOI22_X1 U3137 ( .A1(n3603), .A2(\xmem_inst/mem[10][12] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][12] ), .ZN(n3027) );
  AOI22_X1 U3138 ( .A1(n3585), .A2(\xmem_inst/mem[16][12] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][12] ), .ZN(n3026) );
  NAND4_X1 U3139 ( .A1(n3029), .A2(n3028), .A3(n3027), .A4(n3026), .ZN(n3040)
         );
  AOI22_X1 U3140 ( .A1(n3616), .A2(\xmem_inst/mem[14][12] ), .B1(n3584), .B2(
        \xmem_inst/mem[20][12] ), .ZN(n3033) );
  AOI22_X1 U3141 ( .A1(n3631), .A2(\xmem_inst/mem[34][12] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][12] ), .ZN(n3032) );
  AOI22_X1 U3142 ( .A1(n3624), .A2(\xmem_inst/mem[11][12] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][12] ), .ZN(n3031) );
  AOI22_X1 U3143 ( .A1(n3568), .A2(\xmem_inst/mem[18][12] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][12] ), .ZN(n3030) );
  NAND4_X1 U3144 ( .A1(n3033), .A2(n3032), .A3(n3031), .A4(n3030), .ZN(n3039)
         );
  AOI22_X1 U3145 ( .A1(n3580), .A2(\xmem_inst/mem[38][12] ), .B1(n3613), .B2(
        \xmem_inst/mem[37][12] ), .ZN(n3037) );
  AOI22_X1 U3146 ( .A1(n3626), .A2(\xmem_inst/mem[3][12] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][12] ), .ZN(n3036) );
  AOI22_X1 U3147 ( .A1(n3233), .A2(\xmem_inst/mem[0][12] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][12] ), .ZN(n3035) );
  AOI22_X1 U3148 ( .A1(n3574), .A2(\xmem_inst/mem[27][12] ), .B1(n3629), .B2(
        \xmem_inst/mem[31][12] ), .ZN(n3034) );
  NAND4_X1 U3149 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n3038)
         );
  NOR4_X1 U3150 ( .A1(n3041), .A2(n3040), .A3(n3039), .A4(n3038), .ZN(n3049)
         );
  AOI22_X1 U3151 ( .A1(n3592), .A2(\xmem_inst/mem[41][12] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][12] ), .ZN(n3048) );
  AOI22_X1 U3152 ( .A1(n3627), .A2(\xmem_inst/mem[39][12] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][12] ), .ZN(n3047) );
  AOI22_X1 U3153 ( .A1(n3625), .A2(\xmem_inst/mem[6][12] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][12] ), .ZN(n3045) );
  AOI22_X1 U3154 ( .A1(n3179), .A2(\xmem_inst/mem[8][12] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][12] ), .ZN(n3044) );
  AOI22_X1 U3155 ( .A1(n3252), .A2(\xmem_inst/mem[15][12] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][12] ), .ZN(n3043) );
  AOI22_X1 U3156 ( .A1(n3615), .A2(\xmem_inst/mem[2][12] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][12] ), .ZN(n3042) );
  AND4_X1 U3157 ( .A1(n3045), .A2(n3044), .A3(n3043), .A4(n3042), .ZN(n3046)
         );
  NAND4_X1 U3158 ( .A1(n3049), .A2(n3048), .A3(n3047), .A4(n3046), .ZN(
        \xmem_inst/N267 ) );
  AOI22_X1 U3159 ( .A1(n3597), .A2(\xmem_inst/mem[35][6] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][6] ), .ZN(n3053) );
  AOI22_X1 U3160 ( .A1(n3614), .A2(\xmem_inst/mem[23][6] ), .B1(n3573), .B2(
        \xmem_inst/mem[29][6] ), .ZN(n3052) );
  AOI22_X1 U3161 ( .A1(n3568), .A2(\xmem_inst/mem[18][6] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][6] ), .ZN(n3051) );
  AOI22_X1 U3162 ( .A1(n3631), .A2(\xmem_inst/mem[34][6] ), .B1(n3252), .B2(
        \xmem_inst/mem[15][6] ), .ZN(n3050) );
  NAND4_X1 U3163 ( .A1(n3053), .A2(n3052), .A3(n3051), .A4(n3050), .ZN(n3067)
         );
  AOI22_X1 U3164 ( .A1(n3627), .A2(\xmem_inst/mem[39][6] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][6] ), .ZN(n3057) );
  AOI22_X1 U3165 ( .A1(n3615), .A2(\xmem_inst/mem[2][6] ), .B1(n3574), .B2(
        \xmem_inst/mem[27][6] ), .ZN(n3056) );
  AOI22_X1 U3166 ( .A1(n3598), .A2(\xmem_inst/mem[0][6] ), .B1(n3184), .B2(
        \xmem_inst/mem[37][6] ), .ZN(n3055) );
  AOI22_X1 U3167 ( .A1(n3584), .A2(\xmem_inst/mem[20][6] ), .B1(n3599), .B2(
        \xmem_inst/mem[33][6] ), .ZN(n3054) );
  NAND4_X1 U3168 ( .A1(n3057), .A2(n3056), .A3(n3055), .A4(n3054), .ZN(n3066)
         );
  AOI22_X1 U3169 ( .A1(n3219), .A2(\xmem_inst/mem[9][6] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][6] ), .ZN(n3059) );
  AOI22_X1 U3170 ( .A1(n3593), .A2(\xmem_inst/mem[40][6] ), .B1(n3581), .B2(
        \xmem_inst/mem[22][6] ), .ZN(n3058) );
  NAND2_X1 U3171 ( .A1(n3059), .A2(n3058), .ZN(n3065) );
  AOI22_X1 U3172 ( .A1(n3604), .A2(\xmem_inst/mem[4][6] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][6] ), .ZN(n3063) );
  AOI22_X1 U3173 ( .A1(n3626), .A2(\xmem_inst/mem[3][6] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][6] ), .ZN(n3062) );
  AOI22_X1 U3174 ( .A1(n3585), .A2(\xmem_inst/mem[16][6] ), .B1(n3603), .B2(
        \xmem_inst/mem[10][6] ), .ZN(n3061) );
  AOI22_X1 U3175 ( .A1(n3624), .A2(\xmem_inst/mem[11][6] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][6] ), .ZN(n3060) );
  NAND4_X1 U3176 ( .A1(n3063), .A2(n3062), .A3(n3061), .A4(n3060), .ZN(n3064)
         );
  NOR4_X1 U3177 ( .A1(n3067), .A2(n3066), .A3(n3065), .A4(n3064), .ZN(n3080)
         );
  AOI22_X1 U3178 ( .A1(n3592), .A2(\xmem_inst/mem[41][6] ), .B1(n3220), .B2(
        \xmem_inst/mem[36][6] ), .ZN(n3079) );
  AOI22_X1 U3179 ( .A1(n3253), .A2(\xmem_inst/mem[24][6] ), .B1(n3203), .B2(
        \xmem_inst/mem[38][6] ), .ZN(n3071) );
  NAND2_X1 U3180 ( .A1(n3617), .A2(\xmem_inst/mem[42][6] ), .ZN(n3070) );
  NAND2_X1 U3181 ( .A1(n3616), .A2(\xmem_inst/mem[14][6] ), .ZN(n3069) );
  NAND2_X1 U3182 ( .A1(n3602), .A2(\xmem_inst/mem[32][6] ), .ZN(n3068) );
  AND4_X1 U3183 ( .A1(n3071), .A2(n3070), .A3(n3069), .A4(n3068), .ZN(n3078)
         );
  AOI22_X1 U3184 ( .A1(n3625), .A2(\xmem_inst/mem[6][6] ), .B1(n3072), .B2(
        \xmem_inst/mem[31][6] ), .ZN(n3076) );
  AOI22_X1 U3185 ( .A1(n3571), .A2(\xmem_inst/mem[28][6] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][6] ), .ZN(n3075) );
  AOI22_X1 U3186 ( .A1(n3600), .A2(\xmem_inst/mem[21][6] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][6] ), .ZN(n3074) );
  AOI22_X1 U3187 ( .A1(n3594), .A2(\xmem_inst/mem[19][6] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][6] ), .ZN(n3073) );
  AND4_X1 U3188 ( .A1(n3076), .A2(n3075), .A3(n3074), .A4(n3073), .ZN(n3077)
         );
  NAND4_X1 U3189 ( .A1(n3080), .A2(n3079), .A3(n3078), .A4(n3077), .ZN(
        \xmem_inst/N273 ) );
  NAND2_X1 U3190 ( .A1(n3245), .A2(\xmem_inst/mem[42][8] ), .ZN(n3081) );
  OAI21_X1 U3191 ( .B1(n3082), .B2(n4108), .A(n3081), .ZN(n3083) );
  AOI21_X1 U3192 ( .B1(n3220), .B2(\xmem_inst/mem[36][8] ), .A(n3083), .ZN(
        n3087) );
  AOI22_X1 U3193 ( .A1(n3244), .A2(\xmem_inst/mem[29][8] ), .B1(n3190), .B2(
        \xmem_inst/mem[41][8] ), .ZN(n3086) );
  AOI22_X1 U3194 ( .A1(n3148), .A2(\xmem_inst/mem[32][8] ), .B1(n3084), .B2(
        \xmem_inst/mem[16][8] ), .ZN(n3085) );
  NAND3_X1 U3195 ( .A1(n3087), .A2(n3086), .A3(n3085), .ZN(n3104) );
  AOI22_X1 U3196 ( .A1(n3631), .A2(\xmem_inst/mem[34][8] ), .B1(n3154), .B2(
        \xmem_inst/mem[14][8] ), .ZN(n3091) );
  AOI22_X1 U3197 ( .A1(n3203), .A2(\xmem_inst/mem[38][8] ), .B1(n3153), .B2(
        \xmem_inst/mem[18][8] ), .ZN(n3090) );
  AOI22_X1 U3198 ( .A1(n3254), .A2(\xmem_inst/mem[11][8] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][8] ), .ZN(n3089) );
  AOI22_X1 U3199 ( .A1(n3613), .A2(\xmem_inst/mem[37][8] ), .B1(n3219), .B2(
        \xmem_inst/mem[9][8] ), .ZN(n3088) );
  NAND4_X1 U3200 ( .A1(n3091), .A2(n3090), .A3(n3089), .A4(n3088), .ZN(n3103)
         );
  AOI22_X1 U3201 ( .A1(n3235), .A2(\xmem_inst/mem[6][8] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][8] ), .ZN(n3095) );
  AOI22_X1 U3202 ( .A1(n3600), .A2(\xmem_inst/mem[21][8] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][8] ), .ZN(n3094) );
  AOI22_X1 U3203 ( .A1(n3594), .A2(\xmem_inst/mem[19][8] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][8] ), .ZN(n3093) );
  AOI22_X1 U3204 ( .A1(n3615), .A2(\xmem_inst/mem[2][8] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][8] ), .ZN(n3092) );
  NAND4_X1 U3205 ( .A1(n3095), .A2(n3094), .A3(n3093), .A4(n3092), .ZN(n3102)
         );
  AOI22_X1 U3206 ( .A1(n3598), .A2(\xmem_inst/mem[0][8] ), .B1(n3226), .B2(
        \xmem_inst/mem[33][8] ), .ZN(n3100) );
  AOI22_X1 U3207 ( .A1(n3626), .A2(\xmem_inst/mem[3][8] ), .B1(n3581), .B2(
        \xmem_inst/mem[22][8] ), .ZN(n3099) );
  AOI22_X1 U3208 ( .A1(n3574), .A2(\xmem_inst/mem[27][8] ), .B1(n3096), .B2(
        \xmem_inst/mem[10][8] ), .ZN(n3098) );
  AOI22_X1 U3209 ( .A1(n3252), .A2(\xmem_inst/mem[15][8] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][8] ), .ZN(n3097) );
  NAND4_X1 U3210 ( .A1(n3100), .A2(n3099), .A3(n3098), .A4(n3097), .ZN(n3101)
         );
  NOR4_X1 U3211 ( .A1(n3104), .A2(n3103), .A3(n3102), .A4(n3101), .ZN(n3112)
         );
  AOI22_X1 U3212 ( .A1(n3593), .A2(\xmem_inst/mem[40][8] ), .B1(n3628), .B2(
        \xmem_inst/mem[1][8] ), .ZN(n3111) );
  AOI22_X1 U3213 ( .A1(n3629), .A2(\xmem_inst/mem[31][8] ), .B1(n3253), .B2(
        \xmem_inst/mem[24][8] ), .ZN(n3110) );
  AOI22_X1 U3214 ( .A1(n3614), .A2(\xmem_inst/mem[23][8] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][8] ), .ZN(n3108) );
  AOI22_X1 U3215 ( .A1(n3572), .A2(\xmem_inst/mem[25][8] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][8] ), .ZN(n3107) );
  AOI22_X1 U3216 ( .A1(n3627), .A2(\xmem_inst/mem[39][8] ), .B1(n3251), .B2(
        \xmem_inst/mem[20][8] ), .ZN(n3106) );
  AOI22_X1 U3217 ( .A1(n3597), .A2(\xmem_inst/mem[35][8] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][8] ), .ZN(n3105) );
  AND4_X1 U3218 ( .A1(n3108), .A2(n3107), .A3(n3106), .A4(n3105), .ZN(n3109)
         );
  NAND4_X1 U3219 ( .A1(n3112), .A2(n3111), .A3(n3110), .A4(n3109), .ZN(
        \xmem_inst/N271 ) );
  NAND2_X1 U3220 ( .A1(n3190), .A2(\xmem_inst/mem[41][4] ), .ZN(n3113) );
  OAI21_X1 U3221 ( .B1(n3114), .B2(n4109), .A(n3113), .ZN(n3115) );
  AOI21_X1 U3222 ( .B1(n3193), .B2(\xmem_inst/mem[22][4] ), .A(n3115), .ZN(
        n3118) );
  AOI22_X1 U3223 ( .A1(n3597), .A2(\xmem_inst/mem[35][4] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][4] ), .ZN(n3117) );
  AOI22_X1 U3224 ( .A1(n3630), .A2(\xmem_inst/mem[30][4] ), .B1(n3594), .B2(
        \xmem_inst/mem[19][4] ), .ZN(n3116) );
  NAND3_X1 U3225 ( .A1(n3118), .A2(n3117), .A3(n3116), .ZN(n3134) );
  AOI22_X1 U3226 ( .A1(n3572), .A2(\xmem_inst/mem[25][4] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][4] ), .ZN(n3122) );
  AOI22_X1 U3227 ( .A1(n3614), .A2(\xmem_inst/mem[23][4] ), .B1(n3580), .B2(
        \xmem_inst/mem[38][4] ), .ZN(n3121) );
  AOI22_X1 U3228 ( .A1(n3148), .A2(\xmem_inst/mem[32][4] ), .B1(n3624), .B2(
        \xmem_inst/mem[11][4] ), .ZN(n3120) );
  AOI22_X1 U3229 ( .A1(n3613), .A2(\xmem_inst/mem[37][4] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][4] ), .ZN(n3119) );
  NAND4_X1 U3230 ( .A1(n3122), .A2(n3121), .A3(n3120), .A4(n3119), .ZN(n3133)
         );
  AOI22_X1 U3231 ( .A1(n3629), .A2(\xmem_inst/mem[31][4] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][4] ), .ZN(n3126) );
  AOI22_X1 U3232 ( .A1(n3631), .A2(\xmem_inst/mem[34][4] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][4] ), .ZN(n3125) );
  AOI22_X1 U3233 ( .A1(n3598), .A2(\xmem_inst/mem[0][4] ), .B1(n3628), .B2(
        \xmem_inst/mem[1][4] ), .ZN(n3124) );
  AOI22_X1 U3234 ( .A1(n3252), .A2(\xmem_inst/mem[15][4] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][4] ), .ZN(n3123) );
  NAND4_X1 U3235 ( .A1(n3126), .A2(n3125), .A3(n3124), .A4(n3123), .ZN(n3132)
         );
  AOI22_X1 U3236 ( .A1(n3250), .A2(\xmem_inst/mem[27][4] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][4] ), .ZN(n3130) );
  AOI22_X1 U3237 ( .A1(n3244), .A2(\xmem_inst/mem[29][4] ), .B1(n3619), .B2(
        \xmem_inst/mem[9][4] ), .ZN(n3129) );
  AOI22_X1 U3238 ( .A1(n3253), .A2(\xmem_inst/mem[24][4] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][4] ), .ZN(n3128) );
  AOI22_X1 U3239 ( .A1(n3568), .A2(\xmem_inst/mem[18][4] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][4] ), .ZN(n3127) );
  NAND4_X1 U3240 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .ZN(n3131)
         );
  NOR4_X1 U3241 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n3142)
         );
  AOI22_X1 U3242 ( .A1(n3604), .A2(\xmem_inst/mem[4][4] ), .B1(n3599), .B2(
        \xmem_inst/mem[33][4] ), .ZN(n3141) );
  AOI22_X1 U3243 ( .A1(n3593), .A2(\xmem_inst/mem[40][4] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][4] ), .ZN(n3140) );
  AOI22_X1 U3244 ( .A1(n3615), .A2(\xmem_inst/mem[2][4] ), .B1(n3600), .B2(
        \xmem_inst/mem[21][4] ), .ZN(n3138) );
  AOI22_X1 U3245 ( .A1(n3625), .A2(\xmem_inst/mem[6][4] ), .B1(n3603), .B2(
        \xmem_inst/mem[10][4] ), .ZN(n3137) );
  AOI22_X1 U3246 ( .A1(n3616), .A2(\xmem_inst/mem[14][4] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][4] ), .ZN(n3136) );
  AOI22_X1 U3247 ( .A1(n3584), .A2(\xmem_inst/mem[20][4] ), .B1(n3591), .B2(
        \xmem_inst/mem[8][4] ), .ZN(n3135) );
  AND4_X1 U3248 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3139)
         );
  NAND4_X1 U3249 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(
        \xmem_inst/N275 ) );
  AOI22_X1 U3250 ( .A1(n3626), .A2(\xmem_inst/mem[3][5] ), .B1(n3219), .B2(
        \xmem_inst/mem[9][5] ), .ZN(n3146) );
  AOI22_X1 U3251 ( .A1(n3582), .A2(\xmem_inst/mem[7][5] ), .B1(n3599), .B2(
        \xmem_inst/mem[33][5] ), .ZN(n3145) );
  AOI22_X1 U3252 ( .A1(n3586), .A2(\xmem_inst/mem[24][5] ), .B1(n3603), .B2(
        \xmem_inst/mem[10][5] ), .ZN(n3144) );
  AOI22_X1 U3253 ( .A1(n3625), .A2(\xmem_inst/mem[6][5] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][5] ), .ZN(n3143) );
  NAND4_X1 U3254 ( .A1(n3146), .A2(n3145), .A3(n3144), .A4(n3143), .ZN(n3166)
         );
  AOI22_X1 U3255 ( .A1(n3594), .A2(\xmem_inst/mem[19][5] ), .B1(n3591), .B2(
        \xmem_inst/mem[8][5] ), .ZN(n3152) );
  AOI22_X1 U3256 ( .A1(n3148), .A2(\xmem_inst/mem[32][5] ), .B1(n3147), .B2(
        \xmem_inst/mem[25][5] ), .ZN(n3151) );
  AOI22_X1 U3257 ( .A1(n3598), .A2(\xmem_inst/mem[0][5] ), .B1(n3225), .B2(
        \xmem_inst/mem[5][5] ), .ZN(n3150) );
  AOI22_X1 U3258 ( .A1(n3250), .A2(\xmem_inst/mem[27][5] ), .B1(n3573), .B2(
        \xmem_inst/mem[29][5] ), .ZN(n3149) );
  NAND4_X1 U3259 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3165)
         );
  AOI22_X1 U3260 ( .A1(n3627), .A2(\xmem_inst/mem[39][5] ), .B1(n3153), .B2(
        \xmem_inst/mem[18][5] ), .ZN(n3158) );
  AOI22_X1 U3261 ( .A1(n3615), .A2(\xmem_inst/mem[2][5] ), .B1(n3154), .B2(
        \xmem_inst/mem[14][5] ), .ZN(n3157) );
  AOI22_X1 U3262 ( .A1(n3597), .A2(\xmem_inst/mem[35][5] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][5] ), .ZN(n3156) );
  AOI22_X1 U3263 ( .A1(n3631), .A2(\xmem_inst/mem[34][5] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][5] ), .ZN(n3155) );
  NAND4_X1 U3264 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n3164)
         );
  AOI22_X1 U3265 ( .A1(n3624), .A2(\xmem_inst/mem[11][5] ), .B1(n3604), .B2(
        \xmem_inst/mem[4][5] ), .ZN(n3162) );
  AOI22_X1 U3266 ( .A1(n3614), .A2(\xmem_inst/mem[23][5] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][5] ), .ZN(n3161) );
  AOI22_X1 U3267 ( .A1(n3629), .A2(\xmem_inst/mem[31][5] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][5] ), .ZN(n3160) );
  AOI22_X1 U3268 ( .A1(n3613), .A2(\xmem_inst/mem[37][5] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][5] ), .ZN(n3159) );
  NAND4_X1 U3269 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3163)
         );
  NOR4_X1 U3270 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3176)
         );
  AOI22_X1 U3271 ( .A1(n3580), .A2(\xmem_inst/mem[38][5] ), .B1(n3584), .B2(
        \xmem_inst/mem[20][5] ), .ZN(n3168) );
  AOI22_X1 U3272 ( .A1(n3600), .A2(\xmem_inst/mem[21][5] ), .B1(n3245), .B2(
        \xmem_inst/mem[42][5] ), .ZN(n3167) );
  AND2_X1 U3273 ( .A1(n3168), .A2(n3167), .ZN(n3175) );
  AOI22_X1 U3274 ( .A1(n3592), .A2(\xmem_inst/mem[41][5] ), .B1(n3570), .B2(
        \xmem_inst/mem[17][5] ), .ZN(n3174) );
  AOI22_X1 U3275 ( .A1(n3628), .A2(\xmem_inst/mem[1][5] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][5] ), .ZN(n3172) );
  NAND2_X1 U3276 ( .A1(n3593), .A2(\xmem_inst/mem[40][5] ), .ZN(n3171) );
  NAND2_X1 U3277 ( .A1(n3252), .A2(\xmem_inst/mem[15][5] ), .ZN(n3170) );
  NAND2_X1 U3278 ( .A1(n3220), .A2(\xmem_inst/mem[36][5] ), .ZN(n3169) );
  AND4_X1 U3279 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3173)
         );
  NAND4_X1 U3280 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(
        \xmem_inst/N274 ) );
  AOI22_X1 U3281 ( .A1(n3619), .A2(\xmem_inst/mem[9][0] ), .B1(n3177), .B2(
        \xmem_inst/mem[12][0] ), .ZN(n3183) );
  AOI22_X1 U3282 ( .A1(n3254), .A2(\xmem_inst/mem[11][0] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][0] ), .ZN(n3182) );
  AOI22_X1 U3283 ( .A1(n3600), .A2(\xmem_inst/mem[21][0] ), .B1(n3178), .B2(
        \xmem_inst/mem[30][0] ), .ZN(n3181) );
  AOI22_X1 U3284 ( .A1(n3615), .A2(\xmem_inst/mem[2][0] ), .B1(n3179), .B2(
        \xmem_inst/mem[8][0] ), .ZN(n3180) );
  NAND4_X1 U3285 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3201)
         );
  AOI22_X1 U3286 ( .A1(n3603), .A2(\xmem_inst/mem[10][0] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][0] ), .ZN(n3188) );
  AOI22_X1 U3287 ( .A1(n3626), .A2(\xmem_inst/mem[3][0] ), .B1(n3184), .B2(
        \xmem_inst/mem[37][0] ), .ZN(n3187) );
  AOI22_X1 U3288 ( .A1(n3625), .A2(\xmem_inst/mem[6][0] ), .B1(n3252), .B2(
        \xmem_inst/mem[15][0] ), .ZN(n3186) );
  AOI22_X1 U3289 ( .A1(n3627), .A2(\xmem_inst/mem[39][0] ), .B1(n3251), .B2(
        \xmem_inst/mem[20][0] ), .ZN(n3185) );
  NAND4_X1 U3290 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3200)
         );
  AOI22_X1 U3291 ( .A1(n3245), .A2(\xmem_inst/mem[42][0] ), .B1(n3189), .B2(
        \xmem_inst/mem[28][0] ), .ZN(n3192) );
  AOI22_X1 U3292 ( .A1(n3631), .A2(\xmem_inst/mem[34][0] ), .B1(n3190), .B2(
        \xmem_inst/mem[41][0] ), .ZN(n3191) );
  NAND2_X1 U3293 ( .A1(n3192), .A2(n3191), .ZN(n3199) );
  AOI22_X1 U3294 ( .A1(n3602), .A2(\xmem_inst/mem[32][0] ), .B1(n2295), .B2(
        \xmem_inst/mem[1][0] ), .ZN(n3197) );
  AOI22_X1 U3295 ( .A1(n3598), .A2(\xmem_inst/mem[0][0] ), .B1(n3582), .B2(
        \xmem_inst/mem[7][0] ), .ZN(n3196) );
  AOI22_X1 U3296 ( .A1(n3253), .A2(\xmem_inst/mem[24][0] ), .B1(n3244), .B2(
        \xmem_inst/mem[29][0] ), .ZN(n3195) );
  AOI22_X1 U3297 ( .A1(n3568), .A2(\xmem_inst/mem[18][0] ), .B1(n3193), .B2(
        \xmem_inst/mem[22][0] ), .ZN(n3194) );
  NAND4_X1 U3298 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), .ZN(n3198)
         );
  NOR4_X1 U3299 ( .A1(n3201), .A2(n3200), .A3(n3199), .A4(n3198), .ZN(n3218)
         );
  AOI22_X1 U3300 ( .A1(n3616), .A2(\xmem_inst/mem[14][0] ), .B1(n3202), .B2(
        \xmem_inst/mem[4][0] ), .ZN(n3217) );
  AOI22_X1 U3301 ( .A1(n3572), .A2(\xmem_inst/mem[25][0] ), .B1(n3203), .B2(
        \xmem_inst/mem[38][0] ), .ZN(n3207) );
  NAND2_X1 U3302 ( .A1(n3593), .A2(\xmem_inst/mem[40][0] ), .ZN(n3206) );
  NAND2_X1 U3303 ( .A1(n3574), .A2(\xmem_inst/mem[27][0] ), .ZN(n3205) );
  NAND2_X1 U3304 ( .A1(n3225), .A2(\xmem_inst/mem[5][0] ), .ZN(n3204) );
  AND4_X1 U3305 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3216)
         );
  AOI22_X1 U3306 ( .A1(n3597), .A2(\xmem_inst/mem[35][0] ), .B1(n3208), .B2(
        \xmem_inst/mem[26][0] ), .ZN(n3214) );
  AOI22_X1 U3307 ( .A1(n3629), .A2(\xmem_inst/mem[31][0] ), .B1(n3209), .B2(
        \xmem_inst/mem[17][0] ), .ZN(n3213) );
  AOI22_X1 U3308 ( .A1(n3614), .A2(\xmem_inst/mem[23][0] ), .B1(n3210), .B2(
        \xmem_inst/mem[13][0] ), .ZN(n3212) );
  AOI22_X1 U3309 ( .A1(n3594), .A2(\xmem_inst/mem[19][0] ), .B1(n3599), .B2(
        \xmem_inst/mem[33][0] ), .ZN(n3211) );
  AND4_X1 U3310 ( .A1(n3214), .A2(n3213), .A3(n3212), .A4(n3211), .ZN(n3215)
         );
  NAND4_X1 U3311 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(
        \xmem_inst/N279 ) );
  AOI22_X1 U3312 ( .A1(\xmem_inst/mem[10][31] ), .A2(n3603), .B1(
        \xmem_inst/mem[25][31] ), .B2(n3572), .ZN(n3224) );
  AOI22_X1 U3313 ( .A1(\xmem_inst/mem[1][31] ), .A2(n3628), .B1(
        \xmem_inst/mem[9][31] ), .B2(n3219), .ZN(n3223) );
  AOI22_X1 U3314 ( .A1(\xmem_inst/mem[28][31] ), .A2(n3571), .B1(
        \xmem_inst/mem[30][31] ), .B2(n3630), .ZN(n3222) );
  AOI22_X1 U3315 ( .A1(\xmem_inst/mem[36][31] ), .A2(n3220), .B1(
        \xmem_inst/mem[8][31] ), .B2(n3591), .ZN(n3221) );
  NAND4_X1 U3316 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(n3243)
         );
  AOI22_X1 U3317 ( .A1(\xmem_inst/mem[22][31] ), .A2(n3581), .B1(
        \xmem_inst/mem[17][31] ), .B2(n3570), .ZN(n3230) );
  AOI22_X1 U3318 ( .A1(\xmem_inst/mem[5][31] ), .A2(n3225), .B1(
        \xmem_inst/mem[7][31] ), .B2(n3582), .ZN(n3229) );
  AOI22_X1 U3319 ( .A1(\xmem_inst/mem[33][31] ), .A2(n3226), .B1(
        \xmem_inst/mem[12][31] ), .B2(n3583), .ZN(n3228) );
  AOI22_X1 U3320 ( .A1(\xmem_inst/mem[26][31] ), .A2(n3601), .B1(
        \xmem_inst/mem[13][31] ), .B2(n3569), .ZN(n3227) );
  NAND4_X1 U3321 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3242)
         );
  AOI22_X1 U3322 ( .A1(\xmem_inst/mem[41][31] ), .A2(n3592), .B1(
        \xmem_inst/mem[3][31] ), .B2(n3626), .ZN(n3232) );
  AOI22_X1 U3323 ( .A1(\xmem_inst/mem[4][31] ), .A2(n3604), .B1(
        \xmem_inst/mem[40][31] ), .B2(n3593), .ZN(n3231) );
  NAND2_X1 U3324 ( .A1(n3232), .A2(n3231), .ZN(n3241) );
  AOI22_X1 U3325 ( .A1(\xmem_inst/mem[39][31] ), .A2(n3627), .B1(
        \xmem_inst/mem[34][31] ), .B2(n3631), .ZN(n3239) );
  AOI22_X1 U3326 ( .A1(\xmem_inst/mem[0][31] ), .A2(n3233), .B1(
        \xmem_inst/mem[23][31] ), .B2(n3614), .ZN(n3238) );
  AOI22_X1 U3327 ( .A1(\xmem_inst/mem[6][31] ), .A2(n3235), .B1(
        \xmem_inst/mem[2][31] ), .B2(n3234), .ZN(n3237) );
  AOI22_X1 U3328 ( .A1(\xmem_inst/mem[38][31] ), .A2(n3580), .B1(
        \xmem_inst/mem[35][31] ), .B2(n3597), .ZN(n3236) );
  NAND4_X1 U3329 ( .A1(n3239), .A2(n3238), .A3(n3237), .A4(n3236), .ZN(n3240)
         );
  NOR4_X1 U3330 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3262)
         );
  AOI22_X1 U3331 ( .A1(\xmem_inst/mem[19][31] ), .A2(n3594), .B1(
        \xmem_inst/mem[37][31] ), .B2(n3613), .ZN(n3261) );
  AOI22_X1 U3332 ( .A1(n3244), .A2(\xmem_inst/mem[29][31] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][31] ), .ZN(n3249) );
  NAND2_X1 U3333 ( .A1(\xmem_inst/mem[42][31] ), .A2(n3245), .ZN(n3248) );
  NAND2_X1 U3334 ( .A1(n3568), .A2(\xmem_inst/mem[18][31] ), .ZN(n3247) );
  NAND2_X1 U3335 ( .A1(n3600), .A2(\xmem_inst/mem[21][31] ), .ZN(n3246) );
  AND4_X1 U3336 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3260)
         );
  AOI22_X1 U3337 ( .A1(\xmem_inst/mem[27][31] ), .A2(n3250), .B1(
        \xmem_inst/mem[14][31] ), .B2(n3616), .ZN(n3258) );
  AOI22_X1 U3338 ( .A1(\xmem_inst/mem[15][31] ), .A2(n3252), .B1(
        \xmem_inst/mem[20][31] ), .B2(n3251), .ZN(n3257) );
  AOI22_X1 U3339 ( .A1(\xmem_inst/mem[31][31] ), .A2(n3629), .B1(
        \xmem_inst/mem[32][31] ), .B2(n3602), .ZN(n3256) );
  AOI22_X1 U3340 ( .A1(\xmem_inst/mem[11][31] ), .A2(n3254), .B1(
        \xmem_inst/mem[24][31] ), .B2(n3253), .ZN(n3255) );
  AND4_X1 U3341 ( .A1(n3258), .A2(n3257), .A3(n3256), .A4(n3255), .ZN(n3259)
         );
  NAND4_X1 U3342 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(
        \xmem_inst/N248 ) );
  NAND2_X2 U3343 ( .A1(n3291), .A2(m_valid_y), .ZN(n3537) );
  NOR2_X1 U3344 ( .A1(\mac_unit_inst/adder_reg [2]), .A2(
        \mac_unit_inst/x_mult_f_reg [2]), .ZN(n3518) );
  NOR2_X1 U3345 ( .A1(\mac_unit_inst/adder_reg [3]), .A2(
        \mac_unit_inst/x_mult_f_reg [3]), .ZN(n3520) );
  NOR2_X1 U3346 ( .A1(n3518), .A2(n3520), .ZN(n3264) );
  NOR2_X1 U3347 ( .A1(\mac_unit_inst/adder_reg [1]), .A2(
        \mac_unit_inst/x_mult_f_reg [1]), .ZN(n3530) );
  NAND2_X1 U3348 ( .A1(\mac_unit_inst/adder_reg [0]), .A2(
        \mac_unit_inst/x_mult_f_reg [0]), .ZN(n3533) );
  NAND2_X1 U3349 ( .A1(\mac_unit_inst/adder_reg [1]), .A2(
        \mac_unit_inst/x_mult_f_reg [1]), .ZN(n3531) );
  OAI21_X1 U3350 ( .B1(n3530), .B2(n3533), .A(n3531), .ZN(n3512) );
  NAND2_X1 U3351 ( .A1(\mac_unit_inst/adder_reg [2]), .A2(
        \mac_unit_inst/x_mult_f_reg [2]), .ZN(n3517) );
  NAND2_X1 U3352 ( .A1(\mac_unit_inst/adder_reg [3]), .A2(
        \mac_unit_inst/x_mult_f_reg [3]), .ZN(n3521) );
  OAI21_X1 U3353 ( .B1(n3520), .B2(n3517), .A(n3521), .ZN(n3263) );
  AOI21_X1 U3354 ( .B1(n3264), .B2(n3512), .A(n3263), .ZN(n3366) );
  NOR2_X1 U3355 ( .A1(\mac_unit_inst/adder_reg [4]), .A2(
        \mac_unit_inst/x_mult_f_reg [4]), .ZN(n3489) );
  NOR2_X1 U3356 ( .A1(\mac_unit_inst/adder_reg [5]), .A2(
        \mac_unit_inst/x_mult_f_reg [5]), .ZN(n3498) );
  NOR2_X1 U3357 ( .A1(n3489), .A2(n3498), .ZN(n3368) );
  NOR2_X1 U3358 ( .A1(\mac_unit_inst/adder_reg [6]), .A2(
        \mac_unit_inst/x_mult_f_reg [6]), .ZN(n3505) );
  NOR2_X1 U3359 ( .A1(\mac_unit_inst/adder_reg [7]), .A2(
        \mac_unit_inst/x_mult_f_reg [7]), .ZN(n3369) );
  NOR2_X1 U3360 ( .A1(n3505), .A2(n3369), .ZN(n3266) );
  NAND2_X1 U3361 ( .A1(n3368), .A2(n3266), .ZN(n3268) );
  NAND2_X1 U3362 ( .A1(\mac_unit_inst/adder_reg [4]), .A2(
        \mac_unit_inst/x_mult_f_reg [4]), .ZN(n3494) );
  NAND2_X1 U3363 ( .A1(\mac_unit_inst/adder_reg [5]), .A2(
        \mac_unit_inst/x_mult_f_reg [5]), .ZN(n3499) );
  OAI21_X1 U3364 ( .B1(n3498), .B2(n3494), .A(n3499), .ZN(n3367) );
  NAND2_X1 U3365 ( .A1(\mac_unit_inst/adder_reg [6]), .A2(
        \mac_unit_inst/x_mult_f_reg [6]), .ZN(n3506) );
  NAND2_X1 U3366 ( .A1(\mac_unit_inst/adder_reg [7]), .A2(
        \mac_unit_inst/x_mult_f_reg [7]), .ZN(n3370) );
  OAI21_X1 U3367 ( .B1(n3369), .B2(n3506), .A(n3370), .ZN(n3265) );
  AOI21_X1 U3368 ( .B1(n3266), .B2(n3367), .A(n3265), .ZN(n3267) );
  OAI21_X1 U3369 ( .B1(n3366), .B2(n3268), .A(n3267), .ZN(n3297) );
  NOR2_X1 U3370 ( .A1(\mac_unit_inst/adder_reg [8]), .A2(
        \mac_unit_inst/x_mult_f_reg [8]), .ZN(n3381) );
  NOR2_X1 U3371 ( .A1(\mac_unit_inst/adder_reg [9]), .A2(
        \mac_unit_inst/x_mult_f_reg [9]), .ZN(n3383) );
  NOR2_X1 U3372 ( .A1(n3381), .A2(n3383), .ZN(n3298) );
  NOR2_X1 U3373 ( .A1(\mac_unit_inst/adder_reg [10]), .A2(
        \mac_unit_inst/x_mult_f_reg [10]), .ZN(n3302) );
  NOR2_X1 U3374 ( .A1(\mac_unit_inst/adder_reg [11]), .A2(
        \mac_unit_inst/x_mult_f_reg [11]), .ZN(n3394) );
  NOR2_X1 U3375 ( .A1(n3302), .A2(n3394), .ZN(n3270) );
  NAND2_X1 U3376 ( .A1(n3298), .A2(n3270), .ZN(n3321) );
  NOR2_X1 U3377 ( .A1(\mac_unit_inst/adder_reg [12]), .A2(
        \mac_unit_inst/x_mult_f_reg [12]), .ZN(n3401) );
  NOR2_X1 U3378 ( .A1(\mac_unit_inst/adder_reg [13]), .A2(
        \mac_unit_inst/x_mult_f_reg [13]), .ZN(n3410) );
  NOR2_X1 U3379 ( .A1(n3401), .A2(n3410), .ZN(n3322) );
  NOR2_X1 U3380 ( .A1(\mac_unit_inst/adder_reg [14]), .A2(
        \mac_unit_inst/x_mult_f_reg [14]), .ZN(n3326) );
  NOR2_X1 U3381 ( .A1(\mac_unit_inst/adder_reg [15]), .A2(
        \mac_unit_inst/x_mult_f_reg [15]), .ZN(n3328) );
  NOR2_X1 U3382 ( .A1(n3326), .A2(n3328), .ZN(n3272) );
  NAND2_X1 U3383 ( .A1(n3322), .A2(n3272), .ZN(n3274) );
  NOR2_X1 U3384 ( .A1(n3321), .A2(n3274), .ZN(n3276) );
  NAND2_X1 U3385 ( .A1(\mac_unit_inst/adder_reg [8]), .A2(
        \mac_unit_inst/x_mult_f_reg [8]), .ZN(n3380) );
  NAND2_X1 U3386 ( .A1(\mac_unit_inst/adder_reg [9]), .A2(
        \mac_unit_inst/x_mult_f_reg [9]), .ZN(n3384) );
  OAI21_X1 U3387 ( .B1(n3383), .B2(n3380), .A(n3384), .ZN(n3299) );
  NAND2_X1 U3388 ( .A1(\mac_unit_inst/adder_reg [10]), .A2(
        \mac_unit_inst/x_mult_f_reg [10]), .ZN(n3390) );
  NAND2_X1 U3389 ( .A1(\mac_unit_inst/adder_reg [11]), .A2(
        \mac_unit_inst/x_mult_f_reg [11]), .ZN(n3395) );
  OAI21_X1 U3390 ( .B1(n3394), .B2(n3390), .A(n3395), .ZN(n3269) );
  AOI21_X1 U3391 ( .B1(n3270), .B2(n3299), .A(n3269), .ZN(n3320) );
  NAND2_X1 U3392 ( .A1(\mac_unit_inst/adder_reg [12]), .A2(
        \mac_unit_inst/x_mult_f_reg [12]), .ZN(n3406) );
  NAND2_X1 U3393 ( .A1(\mac_unit_inst/adder_reg [13]), .A2(
        \mac_unit_inst/x_mult_f_reg [13]), .ZN(n3411) );
  OAI21_X1 U3394 ( .B1(n3410), .B2(n3406), .A(n3411), .ZN(n3323) );
  NAND2_X1 U3395 ( .A1(\mac_unit_inst/adder_reg [14]), .A2(
        \mac_unit_inst/x_mult_f_reg [14]), .ZN(n3417) );
  NAND2_X1 U3396 ( .A1(\mac_unit_inst/adder_reg [15]), .A2(
        \mac_unit_inst/x_mult_f_reg [15]), .ZN(n3329) );
  OAI21_X1 U3397 ( .B1(n3328), .B2(n3417), .A(n3329), .ZN(n3271) );
  AOI21_X1 U3398 ( .B1(n3272), .B2(n3323), .A(n3271), .ZN(n3273) );
  OAI21_X1 U3399 ( .B1(n3320), .B2(n3274), .A(n3273), .ZN(n3275) );
  AOI21_X1 U3400 ( .B1(n3297), .B2(n3276), .A(n3275), .ZN(n3335) );
  NOR2_X1 U3401 ( .A1(\mac_unit_inst/adder_reg [16]), .A2(
        \mac_unit_inst/x_mult_f_reg [16]), .ZN(n3336) );
  NOR2_X1 U3402 ( .A1(\mac_unit_inst/adder_reg [17]), .A2(
        \mac_unit_inst/x_mult_f_reg [17]), .ZN(n3343) );
  NOR2_X1 U3403 ( .A1(n3336), .A2(n3343), .ZN(n3351) );
  NOR2_X1 U3404 ( .A1(\mac_unit_inst/adder_reg [18]), .A2(
        \mac_unit_inst/x_mult_f_reg [18]), .ZN(n3357) );
  NOR2_X1 U3405 ( .A1(\mac_unit_inst/adder_reg [19]), .A2(
        \mac_unit_inst/x_mult_f_reg [19]), .ZN(n3359) );
  NOR2_X1 U3406 ( .A1(n3357), .A2(n3359), .ZN(n3278) );
  NAND2_X1 U3407 ( .A1(n3351), .A2(n3278), .ZN(n3424) );
  NOR2_X1 U3408 ( .A1(\mac_unit_inst/adder_reg [20]), .A2(
        \mac_unit_inst/x_mult_f_reg [20]), .ZN(n3433) );
  NOR2_X1 U3409 ( .A1(\mac_unit_inst/adder_reg [21]), .A2(
        \mac_unit_inst/x_mult_f_reg [21]), .ZN(n3435) );
  NOR2_X1 U3410 ( .A1(n3433), .A2(n3435), .ZN(n3443) );
  NOR2_X1 U3411 ( .A1(\mac_unit_inst/adder_reg [22]), .A2(
        \mac_unit_inst/x_mult_f_reg [22]), .ZN(n3450) );
  NOR2_X1 U3412 ( .A1(\mac_unit_inst/adder_reg [23]), .A2(
        \mac_unit_inst/x_mult_f_reg [23]), .ZN(n3452) );
  NOR2_X1 U3413 ( .A1(n3450), .A2(n3452), .ZN(n3280) );
  NAND2_X1 U3414 ( .A1(n3443), .A2(n3280), .ZN(n3282) );
  NOR2_X1 U3415 ( .A1(n3424), .A2(n3282), .ZN(n3460) );
  NOR2_X1 U3416 ( .A1(\mac_unit_inst/adder_reg [24]), .A2(
        \mac_unit_inst/x_mult_f_reg [24]), .ZN(n3467) );
  INV_X1 U3417 ( .A(n3467), .ZN(n3462) );
  NAND2_X1 U3418 ( .A1(n3462), .A2(n3470), .ZN(n3475) );
  NOR2_X1 U3419 ( .A1(\mac_unit_inst/adder_reg [26]), .A2(
        \mac_unit_inst/x_mult_f_reg [26]), .ZN(n3480) );
  NOR2_X1 U3420 ( .A1(n3475), .A2(n3480), .ZN(n3286) );
  NAND2_X1 U3421 ( .A1(n3460), .A2(n3286), .ZN(n3288) );
  NAND2_X1 U3422 ( .A1(\mac_unit_inst/adder_reg [16]), .A2(
        \mac_unit_inst/x_mult_f_reg [16]), .ZN(n3340) );
  NAND2_X1 U3423 ( .A1(\mac_unit_inst/adder_reg [17]), .A2(
        \mac_unit_inst/x_mult_f_reg [17]), .ZN(n3344) );
  OAI21_X1 U3424 ( .B1(n3343), .B2(n3340), .A(n3344), .ZN(n3350) );
  NAND2_X1 U3425 ( .A1(\mac_unit_inst/adder_reg [18]), .A2(
        \mac_unit_inst/x_mult_f_reg [18]), .ZN(n3356) );
  NAND2_X1 U3426 ( .A1(\mac_unit_inst/adder_reg [19]), .A2(
        \mac_unit_inst/x_mult_f_reg [19]), .ZN(n3360) );
  OAI21_X1 U3427 ( .B1(n3359), .B2(n3356), .A(n3360), .ZN(n3277) );
  AOI21_X1 U3428 ( .B1(n3278), .B2(n3350), .A(n3277), .ZN(n3425) );
  NAND2_X1 U3429 ( .A1(\mac_unit_inst/adder_reg [20]), .A2(
        \mac_unit_inst/x_mult_f_reg [20]), .ZN(n3432) );
  NAND2_X1 U3430 ( .A1(\mac_unit_inst/adder_reg [21]), .A2(
        \mac_unit_inst/x_mult_f_reg [21]), .ZN(n3436) );
  OAI21_X1 U3431 ( .B1(n3435), .B2(n3432), .A(n3436), .ZN(n3442) );
  NAND2_X1 U3432 ( .A1(\mac_unit_inst/adder_reg [22]), .A2(
        \mac_unit_inst/x_mult_f_reg [22]), .ZN(n3449) );
  NAND2_X1 U3433 ( .A1(\mac_unit_inst/adder_reg [23]), .A2(
        \mac_unit_inst/x_mult_f_reg [23]), .ZN(n3453) );
  OAI21_X1 U3434 ( .B1(n3452), .B2(n3449), .A(n3453), .ZN(n3279) );
  AOI21_X1 U3435 ( .B1(n3280), .B2(n3442), .A(n3279), .ZN(n3281) );
  OAI21_X1 U3436 ( .B1(n3425), .B2(n3282), .A(n3281), .ZN(n3459) );
  NAND2_X1 U3437 ( .A1(\mac_unit_inst/adder_reg [24]), .A2(
        \mac_unit_inst/x_mult_f_reg [24]), .ZN(n3466) );
  INV_X1 U3438 ( .A(n3466), .ZN(n3284) );
  NAND2_X1 U3439 ( .A1(\mac_unit_inst/adder_reg [25]), .A2(
        \mac_unit_inst/x_mult_f_reg [25]), .ZN(n3469) );
  INV_X1 U3440 ( .A(n3469), .ZN(n3283) );
  AOI21_X1 U3441 ( .B1(n3470), .B2(n3284), .A(n3283), .ZN(n3476) );
  NAND2_X1 U3442 ( .A1(\mac_unit_inst/adder_reg [26]), .A2(
        \mac_unit_inst/x_mult_f_reg [26]), .ZN(n3481) );
  OAI21_X1 U3443 ( .B1(n3476), .B2(n3480), .A(n3481), .ZN(n3285) );
  AOI21_X1 U3444 ( .B1(n3459), .B2(n3286), .A(n3285), .ZN(n3287) );
  OAI21_X1 U3445 ( .B1(n3335), .B2(n3288), .A(n3287), .ZN(n3308) );
  FA_X1 U3446 ( .A(n309), .B(n4112), .CI(n3289), .CO(n3290), .S(n3293) );
  NOR2_X1 U3447 ( .A1(n3293), .A2(n3290), .ZN(n3296) );
  INV_X1 U3448 ( .A(n3306), .ZN(n3292) );
  AND2_X1 U3449 ( .A1(n3291), .A2(n4073), .ZN(n3305) );
  OAI211_X1 U3450 ( .C1(n3296), .C2(n3293), .A(n3292), .B(n3305), .ZN(n3294)
         );
  OAI21_X1 U3451 ( .B1(n309), .B2(n3537), .A(n3294), .ZN(\mac_unit_inst/n81 )
         );
  INV_X1 U3452 ( .A(n3305), .ZN(n3295) );
  INV_X1 U3453 ( .A(n3297), .ZN(n3382) );
  INV_X1 U3454 ( .A(n3298), .ZN(n3301) );
  INV_X1 U3455 ( .A(n3299), .ZN(n3300) );
  OAI21_X1 U3456 ( .B1(n3382), .B2(n3301), .A(n3300), .ZN(n3393) );
  INV_X1 U3457 ( .A(n3302), .ZN(n3392) );
  NAND2_X1 U3458 ( .A1(n3392), .A2(n3390), .ZN(n3303) );
  XNOR2_X1 U3459 ( .A(n3393), .B(n3303), .ZN(n3304) );
  NAND2_X1 U3460 ( .A1(n3422), .A2(n3304), .ZN(n3307) );
  OAI211_X1 U3461 ( .C1(n3537), .C2(n322), .A(n3307), .B(n3492), .ZN(
        \mac_unit_inst/n102 ) );
  FA_X1 U3462 ( .A(\mac_unit_inst/adder_reg [27]), .B(
        \mac_unit_inst/x_mult_f_reg [27]), .CI(n3308), .CO(n3311), .S(n3309)
         );
  NAND2_X1 U3463 ( .A1(n3486), .A2(n3309), .ZN(n3310) );
  OAI211_X1 U3464 ( .C1(n3537), .C2(n318), .A(n3310), .B(n3492), .ZN(
        \mac_unit_inst/n85 ) );
  FA_X1 U3465 ( .A(\mac_unit_inst/adder_reg [28]), .B(
        \mac_unit_inst/x_mult_f_reg [28]), .CI(n3311), .CO(n3314), .S(n3312)
         );
  NAND2_X1 U3466 ( .A1(n3486), .A2(n3312), .ZN(n3313) );
  OAI211_X1 U3467 ( .C1(n3537), .C2(n319), .A(n3313), .B(n3492), .ZN(
        \mac_unit_inst/n84 ) );
  FA_X1 U3468 ( .A(\mac_unit_inst/adder_reg [29]), .B(
        \mac_unit_inst/x_mult_f_reg [29]), .CI(n3314), .CO(n3317), .S(n3315)
         );
  NAND2_X1 U3469 ( .A1(n3486), .A2(n3315), .ZN(n3316) );
  OAI211_X1 U3470 ( .C1(n3537), .C2(n320), .A(n3316), .B(n3492), .ZN(
        \mac_unit_inst/n83 ) );
  FA_X1 U3471 ( .A(\mac_unit_inst/adder_reg [30]), .B(
        \mac_unit_inst/x_mult_f_reg [30]), .CI(n3317), .CO(n3289), .S(n3318)
         );
  NAND2_X1 U3472 ( .A1(n3486), .A2(n3318), .ZN(n3319) );
  OAI211_X1 U3473 ( .C1(n3537), .C2(n321), .A(n3319), .B(n3492), .ZN(
        \mac_unit_inst/n82 ) );
  OAI21_X1 U3474 ( .B1(n3382), .B2(n3321), .A(n3320), .ZN(n3409) );
  INV_X1 U3475 ( .A(n3409), .ZN(n3403) );
  INV_X1 U3476 ( .A(n3322), .ZN(n3325) );
  INV_X1 U3477 ( .A(n3323), .ZN(n3324) );
  OAI21_X1 U3478 ( .B1(n3403), .B2(n3325), .A(n3324), .ZN(n3420) );
  INV_X1 U3479 ( .A(n3326), .ZN(n3418) );
  INV_X1 U3480 ( .A(n3417), .ZN(n3327) );
  AOI21_X1 U3481 ( .B1(n3420), .B2(n3418), .A(n3327), .ZN(n3332) );
  INV_X1 U3482 ( .A(n3328), .ZN(n3330) );
  NAND2_X1 U3483 ( .A1(n3330), .A2(n3329), .ZN(n3331) );
  XOR2_X1 U3484 ( .A(n3332), .B(n3331), .Z(n3333) );
  NAND2_X1 U3485 ( .A1(n3422), .A2(n3333), .ZN(n3334) );
  OAI211_X1 U3486 ( .C1(n3537), .C2(n4093), .A(n3334), .B(n3492), .ZN(
        \mac_unit_inst/n97 ) );
  INV_X1 U3487 ( .A(n3335), .ZN(n3461) );
  INV_X1 U3488 ( .A(n3336), .ZN(n3342) );
  NAND2_X1 U3489 ( .A1(n3342), .A2(n3340), .ZN(n3337) );
  XNOR2_X1 U3490 ( .A(n3461), .B(n3337), .ZN(n3338) );
  NAND2_X1 U3491 ( .A1(n3422), .A2(n3338), .ZN(n3339) );
  OAI211_X1 U3492 ( .C1(n3537), .C2(n4094), .A(n3339), .B(n3492), .ZN(
        \mac_unit_inst/n96 ) );
  INV_X1 U3493 ( .A(n3340), .ZN(n3341) );
  AOI21_X1 U3494 ( .B1(n3461), .B2(n3342), .A(n3341), .ZN(n3347) );
  INV_X1 U3495 ( .A(n3343), .ZN(n3345) );
  NAND2_X1 U3496 ( .A1(n3345), .A2(n3344), .ZN(n3346) );
  XOR2_X1 U3497 ( .A(n3347), .B(n3346), .Z(n3348) );
  NAND2_X1 U3498 ( .A1(n3422), .A2(n3348), .ZN(n3349) );
  OAI211_X1 U3499 ( .C1(n3537), .C2(n4095), .A(n3349), .B(n3492), .ZN(
        \mac_unit_inst/n95 ) );
  AOI21_X1 U3500 ( .B1(n3461), .B2(n3351), .A(n3350), .ZN(n3358) );
  INV_X1 U3501 ( .A(n3357), .ZN(n3352) );
  NAND2_X1 U3502 ( .A1(n3352), .A2(n3356), .ZN(n3353) );
  XOR2_X1 U3503 ( .A(n3358), .B(n3353), .Z(n3354) );
  NAND2_X1 U3504 ( .A1(n3422), .A2(n3354), .ZN(n3355) );
  OAI211_X1 U3505 ( .C1(n3537), .C2(n4096), .A(n3355), .B(n3492), .ZN(
        \mac_unit_inst/n94 ) );
  OAI21_X1 U3506 ( .B1(n3358), .B2(n3357), .A(n3356), .ZN(n3363) );
  INV_X1 U3507 ( .A(n3359), .ZN(n3361) );
  NAND2_X1 U3508 ( .A1(n3361), .A2(n3360), .ZN(n3362) );
  XNOR2_X1 U3509 ( .A(n3363), .B(n3362), .ZN(n3364) );
  NAND2_X1 U3510 ( .A1(n3486), .A2(n3364), .ZN(n3365) );
  OAI211_X1 U3511 ( .C1(n3537), .C2(n4097), .A(n3365), .B(n3492), .ZN(
        \mac_unit_inst/n93 ) );
  INV_X1 U3512 ( .A(n3366), .ZN(n3497) );
  AOI21_X1 U3513 ( .B1(n3497), .B2(n3368), .A(n3367), .ZN(n3509) );
  OAI21_X1 U3514 ( .B1(n3509), .B2(n3505), .A(n3506), .ZN(n3373) );
  INV_X1 U3515 ( .A(n3369), .ZN(n3371) );
  NAND2_X1 U3516 ( .A1(n3371), .A2(n3370), .ZN(n3372) );
  XNOR2_X1 U3517 ( .A(n3373), .B(n3372), .ZN(n3374) );
  NAND2_X1 U3518 ( .A1(n3422), .A2(n3374), .ZN(n3375) );
  OAI211_X1 U3519 ( .C1(n3537), .C2(n4089), .A(n3375), .B(n3492), .ZN(
        \mac_unit_inst/n105 ) );
  INV_X1 U3520 ( .A(n3381), .ZN(n3376) );
  NAND2_X1 U3521 ( .A1(n3376), .A2(n3380), .ZN(n3377) );
  XOR2_X1 U3522 ( .A(n3382), .B(n3377), .Z(n3378) );
  NAND2_X1 U3523 ( .A1(n3422), .A2(n3378), .ZN(n3379) );
  OAI211_X1 U3524 ( .C1(n3537), .C2(n323), .A(n3379), .B(n3492), .ZN(
        \mac_unit_inst/n104 ) );
  OAI21_X1 U3525 ( .B1(n3382), .B2(n3381), .A(n3380), .ZN(n3387) );
  INV_X1 U3526 ( .A(n3383), .ZN(n3385) );
  NAND2_X1 U3527 ( .A1(n3385), .A2(n3384), .ZN(n3386) );
  XNOR2_X1 U3528 ( .A(n3387), .B(n3386), .ZN(n3388) );
  NAND2_X1 U3529 ( .A1(n3422), .A2(n3388), .ZN(n3389) );
  OAI211_X1 U3530 ( .C1(n3537), .C2(n324), .A(n3389), .B(n3492), .ZN(
        \mac_unit_inst/n103 ) );
  INV_X1 U3531 ( .A(n3390), .ZN(n3391) );
  AOI21_X1 U3532 ( .B1(n3393), .B2(n3392), .A(n3391), .ZN(n3398) );
  INV_X1 U3533 ( .A(n3394), .ZN(n3396) );
  NAND2_X1 U3534 ( .A1(n3396), .A2(n3395), .ZN(n3397) );
  XOR2_X1 U3535 ( .A(n3398), .B(n3397), .Z(n3399) );
  NAND2_X1 U3536 ( .A1(n3422), .A2(n3399), .ZN(n3400) );
  OAI211_X1 U3537 ( .C1(n3537), .C2(n325), .A(n3400), .B(n3492), .ZN(
        \mac_unit_inst/n101 ) );
  INV_X1 U3538 ( .A(n3401), .ZN(n3408) );
  NAND2_X1 U3539 ( .A1(n3408), .A2(n3406), .ZN(n3402) );
  XOR2_X1 U3540 ( .A(n3403), .B(n3402), .Z(n3404) );
  NAND2_X1 U3541 ( .A1(n3422), .A2(n3404), .ZN(n3405) );
  OAI211_X1 U3542 ( .C1(n3537), .C2(n4090), .A(n3405), .B(n3492), .ZN(
        \mac_unit_inst/n100 ) );
  INV_X1 U3543 ( .A(n3406), .ZN(n3407) );
  AOI21_X1 U3544 ( .B1(n3409), .B2(n3408), .A(n3407), .ZN(n3414) );
  INV_X1 U3545 ( .A(n3410), .ZN(n3412) );
  NAND2_X1 U3546 ( .A1(n3412), .A2(n3411), .ZN(n3413) );
  XOR2_X1 U3547 ( .A(n3414), .B(n3413), .Z(n3415) );
  NAND2_X1 U3548 ( .A1(n3422), .A2(n3415), .ZN(n3416) );
  OAI211_X1 U3549 ( .C1(n3537), .C2(n4091), .A(n3416), .B(n3492), .ZN(
        \mac_unit_inst/n99 ) );
  NAND2_X1 U3550 ( .A1(n3418), .A2(n3417), .ZN(n3419) );
  XNOR2_X1 U3551 ( .A(n3420), .B(n3419), .ZN(n3421) );
  NAND2_X1 U3552 ( .A1(n3422), .A2(n3421), .ZN(n3423) );
  OAI211_X1 U3553 ( .C1(n3537), .C2(n4092), .A(n3423), .B(n3492), .ZN(
        \mac_unit_inst/n98 ) );
  INV_X1 U3554 ( .A(n3424), .ZN(n3427) );
  INV_X1 U3555 ( .A(n3425), .ZN(n3426) );
  AOI21_X1 U3556 ( .B1(n3461), .B2(n3427), .A(n3426), .ZN(n3434) );
  INV_X1 U3557 ( .A(n3434), .ZN(n3444) );
  INV_X1 U3558 ( .A(n3433), .ZN(n3428) );
  NAND2_X1 U3559 ( .A1(n3428), .A2(n3432), .ZN(n3429) );
  XNOR2_X1 U3560 ( .A(n3444), .B(n3429), .ZN(n3430) );
  NAND2_X1 U3561 ( .A1(n3486), .A2(n3430), .ZN(n3431) );
  OAI211_X1 U3562 ( .C1(n3537), .C2(n4098), .A(n3431), .B(n3492), .ZN(
        \mac_unit_inst/n92 ) );
  OAI21_X1 U3563 ( .B1(n3434), .B2(n3433), .A(n3432), .ZN(n3439) );
  INV_X1 U3564 ( .A(n3435), .ZN(n3437) );
  NAND2_X1 U3565 ( .A1(n3437), .A2(n3436), .ZN(n3438) );
  XNOR2_X1 U3566 ( .A(n3439), .B(n3438), .ZN(n3440) );
  NAND2_X1 U3567 ( .A1(n3486), .A2(n3440), .ZN(n3441) );
  OAI211_X1 U3568 ( .C1(n3537), .C2(n4099), .A(n3441), .B(n3492), .ZN(
        \mac_unit_inst/n91 ) );
  AOI21_X1 U3569 ( .B1(n3444), .B2(n3443), .A(n3442), .ZN(n3451) );
  INV_X1 U3570 ( .A(n3450), .ZN(n3445) );
  NAND2_X1 U3571 ( .A1(n3445), .A2(n3449), .ZN(n3446) );
  XOR2_X1 U3572 ( .A(n3451), .B(n3446), .Z(n3447) );
  NAND2_X1 U3573 ( .A1(n3486), .A2(n3447), .ZN(n3448) );
  OAI211_X1 U3574 ( .C1(n3537), .C2(n4100), .A(n3448), .B(n3492), .ZN(
        \mac_unit_inst/n90 ) );
  OAI21_X1 U3575 ( .B1(n3451), .B2(n3450), .A(n3449), .ZN(n3456) );
  INV_X1 U3576 ( .A(n3452), .ZN(n3454) );
  NAND2_X1 U3577 ( .A1(n3454), .A2(n3453), .ZN(n3455) );
  XNOR2_X1 U3578 ( .A(n3456), .B(n3455), .ZN(n3457) );
  NAND2_X1 U3579 ( .A1(n3486), .A2(n3457), .ZN(n3458) );
  OAI211_X1 U3580 ( .C1(n3537), .C2(n4101), .A(n3458), .B(n3492), .ZN(
        \mac_unit_inst/n89 ) );
  AOI21_X1 U3581 ( .B1(n3461), .B2(n3460), .A(n3459), .ZN(n3468) );
  INV_X1 U3582 ( .A(n3468), .ZN(n3479) );
  NAND2_X1 U3583 ( .A1(n3462), .A2(n3466), .ZN(n3463) );
  XNOR2_X1 U3584 ( .A(n3479), .B(n3463), .ZN(n3464) );
  NAND2_X1 U3585 ( .A1(n3486), .A2(n3464), .ZN(n3465) );
  OAI211_X1 U3586 ( .C1(n3537), .C2(n326), .A(n3465), .B(n3492), .ZN(
        \mac_unit_inst/n88 ) );
  OAI21_X1 U3587 ( .B1(n3468), .B2(n3467), .A(n3466), .ZN(n3472) );
  NAND2_X1 U3588 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  XNOR2_X1 U3589 ( .A(n3472), .B(n3471), .ZN(n3473) );
  NAND2_X1 U3590 ( .A1(n3486), .A2(n3473), .ZN(n3474) );
  OAI211_X1 U3591 ( .C1(n3537), .C2(n327), .A(n3474), .B(n3492), .ZN(
        \mac_unit_inst/n87 ) );
  INV_X1 U3592 ( .A(n3475), .ZN(n3478) );
  INV_X1 U3593 ( .A(n3476), .ZN(n3477) );
  AOI21_X1 U3594 ( .B1(n3479), .B2(n3478), .A(n3477), .ZN(n3484) );
  INV_X1 U3595 ( .A(n3480), .ZN(n3482) );
  NAND2_X1 U3596 ( .A1(n3482), .A2(n3481), .ZN(n3483) );
  XOR2_X1 U3597 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND2_X1 U3598 ( .A1(n3486), .A2(n3485), .ZN(n3487) );
  OAI211_X1 U3599 ( .C1(n3537), .C2(n328), .A(n3487), .B(n3492), .ZN(
        \mac_unit_inst/n86 ) );
  INV_X1 U3600 ( .A(n3489), .ZN(n3496) );
  NAND2_X1 U3601 ( .A1(n3496), .A2(n3494), .ZN(n3490) );
  XNOR2_X1 U3602 ( .A(n3497), .B(n3490), .ZN(n3491) );
  NAND2_X1 U3603 ( .A1(n3488), .A2(n3491), .ZN(n3493) );
  OAI211_X1 U3604 ( .C1(n3537), .C2(n4103), .A(n3493), .B(n3492), .ZN(
        \mac_unit_inst/n108 ) );
  INV_X1 U3605 ( .A(n3494), .ZN(n3495) );
  AOI21_X1 U3606 ( .B1(n3497), .B2(n3496), .A(n3495), .ZN(n3502) );
  INV_X1 U3607 ( .A(n3498), .ZN(n3500) );
  NAND2_X1 U3608 ( .A1(n3500), .A2(n3499), .ZN(n3501) );
  XOR2_X1 U3609 ( .A(n3502), .B(n3501), .Z(n3503) );
  NAND2_X1 U3610 ( .A1(n3422), .A2(n3503), .ZN(n3504) );
  OAI211_X1 U3611 ( .C1(n3537), .C2(n4104), .A(n3504), .B(n3492), .ZN(
        \mac_unit_inst/n107 ) );
  INV_X1 U3612 ( .A(n3505), .ZN(n3507) );
  NAND2_X1 U3613 ( .A1(n3507), .A2(n3506), .ZN(n3508) );
  XOR2_X1 U3614 ( .A(n3509), .B(n3508), .Z(n3510) );
  NAND2_X1 U3615 ( .A1(n3486), .A2(n3510), .ZN(n3511) );
  OAI211_X1 U3616 ( .C1(n3537), .C2(n4088), .A(n3511), .B(n3492), .ZN(
        \mac_unit_inst/n106 ) );
  INV_X1 U3617 ( .A(n3512), .ZN(n3519) );
  INV_X1 U3618 ( .A(n3518), .ZN(n3513) );
  NAND2_X1 U3619 ( .A1(n3513), .A2(n3517), .ZN(n3514) );
  XOR2_X1 U3620 ( .A(n3519), .B(n3514), .Z(n3515) );
  NAND2_X1 U3621 ( .A1(n3488), .A2(n3515), .ZN(n3516) );
  OAI211_X1 U3622 ( .C1(n3537), .C2(n4086), .A(n3516), .B(n3492), .ZN(
        \mac_unit_inst/n110 ) );
  OAI21_X1 U3623 ( .B1(n3519), .B2(n3518), .A(n3517), .ZN(n3524) );
  INV_X1 U3624 ( .A(n3520), .ZN(n3522) );
  NAND2_X1 U3625 ( .A1(n3522), .A2(n3521), .ZN(n3523) );
  XNOR2_X1 U3626 ( .A(n3524), .B(n3523), .ZN(n3525) );
  NAND2_X1 U3627 ( .A1(n3488), .A2(n3525), .ZN(n3526) );
  OAI211_X1 U3628 ( .C1(n3537), .C2(n4087), .A(n3526), .B(n3492), .ZN(
        \mac_unit_inst/n109 ) );
  OR2_X1 U3629 ( .A1(\mac_unit_inst/adder_reg [0]), .A2(
        \mac_unit_inst/x_mult_f_reg [0]), .ZN(n3527) );
  AND2_X1 U3630 ( .A1(n3527), .A2(n3533), .ZN(n3528) );
  NAND2_X1 U3631 ( .A1(n3488), .A2(n3528), .ZN(n3529) );
  OAI211_X1 U3632 ( .C1(n3537), .C2(n4084), .A(n3529), .B(n3492), .ZN(
        \mac_unit_inst/n112 ) );
  INV_X1 U3633 ( .A(n3530), .ZN(n3532) );
  NAND2_X1 U3634 ( .A1(n3532), .A2(n3531), .ZN(n3534) );
  XOR2_X1 U3635 ( .A(n3534), .B(n3533), .Z(n3535) );
  NAND2_X1 U3636 ( .A1(n3488), .A2(n3535), .ZN(n3536) );
  OAI211_X1 U3637 ( .C1(n3537), .C2(n4085), .A(n3536), .B(n3492), .ZN(
        \mac_unit_inst/n111 ) );
  NAND3_X1 U3638 ( .A1(n4075), .A2(n4025), .A3(
        \ctrl_conv_output_inst/m_pre_pre_valid_y ), .ZN(n4013) );
  NAND3_X1 U3639 ( .A1(\ctrl_conv_output_inst/cnt_conv [2]), .A2(
        \ctrl_conv_output_inst/cnt_conv [1]), .A3(
        \ctrl_conv_output_inst/cnt_conv [0]), .ZN(n3540) );
  NOR2_X1 U3640 ( .A1(n4013), .A2(n3540), .ZN(n3539) );
  NAND2_X1 U3641 ( .A1(\ctrl_conv_output_inst/m_pre_pre_valid_y ), .A2(n4075), 
        .ZN(n4015) );
  OAI21_X1 U3642 ( .B1(n4015), .B2(n3540), .A(n4025), .ZN(n3541) );
  INV_X1 U3643 ( .A(n3541), .ZN(n3538) );
  MUX2_X1 U3644 ( .A(n3539), .B(n3538), .S(\ctrl_conv_output_inst/cnt_conv [3]), .Z(n116) );
  OR3_X1 U3645 ( .A1(n4110), .A2(n4013), .A3(n3540), .ZN(n4021) );
  NOR2_X1 U3646 ( .A1(n4076), .A2(n4021), .ZN(n3544) );
  INV_X1 U3647 ( .A(n4013), .ZN(n4016) );
  OAI21_X1 U3648 ( .B1(\ctrl_conv_output_inst/cnt_conv [3]), .B2(n4013), .A(
        n3541), .ZN(n4020) );
  AOI21_X1 U3649 ( .B1(n4016), .B2(n4076), .A(n4020), .ZN(n3542) );
  INV_X1 U3650 ( .A(n3542), .ZN(n3543) );
  MUX2_X1 U3651 ( .A(n3544), .B(n3543), .S(\ctrl_conv_output_inst/cnt_conv [5]), .Z(n120) );
  NAND2_X1 U3652 ( .A1(n3549), .A2(n3545), .ZN(n3551) );
  NOR2_X1 U3653 ( .A1(n3546), .A2(n3551), .ZN(n3554) );
  AOI21_X1 U3654 ( .B1(n3549), .B2(n3548), .A(n3547), .ZN(n3550) );
  OAI21_X1 U3655 ( .B1(n3552), .B2(n3551), .A(n3550), .ZN(n3553) );
  AOI21_X1 U3656 ( .B1(n3554), .B2(n302), .A(n3553), .ZN(n3560) );
  OR2_X1 U3657 ( .A1(n3556), .A2(n3555), .ZN(n3558) );
  NAND2_X1 U3658 ( .A1(n3556), .A2(n3555), .ZN(n3557) );
  NAND2_X1 U3659 ( .A1(n3558), .A2(n3557), .ZN(n3559) );
  XOR2_X1 U3660 ( .A(n3560), .B(n3559), .Z(n3564) );
  INV_X1 U3661 ( .A(n292), .ZN(n3563) );
  OAI211_X1 U3662 ( .C1(n304), .C2(n3564), .A(n3563), .B(n3562), .ZN(n3566) );
  OAI21_X1 U3663 ( .B1(n4112), .B2(n2223), .A(n3566), .ZN(\mac_unit_inst/n144 ) );
  AOI22_X1 U3664 ( .A1(n3568), .A2(\xmem_inst/mem[18][1] ), .B1(n3567), .B2(
        \xmem_inst/mem[5][1] ), .ZN(n3578) );
  AOI22_X1 U3665 ( .A1(n3570), .A2(\xmem_inst/mem[17][1] ), .B1(n3569), .B2(
        \xmem_inst/mem[13][1] ), .ZN(n3577) );
  AOI22_X1 U3666 ( .A1(n3572), .A2(\xmem_inst/mem[25][1] ), .B1(n3571), .B2(
        \xmem_inst/mem[28][1] ), .ZN(n3576) );
  AOI22_X1 U3667 ( .A1(n3574), .A2(\xmem_inst/mem[27][1] ), .B1(n3573), .B2(
        \xmem_inst/mem[29][1] ), .ZN(n3575) );
  NAND4_X1 U3668 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(n3612)
         );
  AOI22_X1 U3669 ( .A1(n3580), .A2(\xmem_inst/mem[38][1] ), .B1(n3579), .B2(
        \xmem_inst/mem[36][1] ), .ZN(n3590) );
  AOI22_X1 U3670 ( .A1(n3582), .A2(\xmem_inst/mem[7][1] ), .B1(n3581), .B2(
        \xmem_inst/mem[22][1] ), .ZN(n3589) );
  AOI22_X1 U3671 ( .A1(n3584), .A2(\xmem_inst/mem[20][1] ), .B1(n3583), .B2(
        \xmem_inst/mem[12][1] ), .ZN(n3588) );
  AOI22_X1 U3672 ( .A1(n3586), .A2(\xmem_inst/mem[24][1] ), .B1(n3585), .B2(
        \xmem_inst/mem[16][1] ), .ZN(n3587) );
  NAND4_X1 U3673 ( .A1(n3590), .A2(n3589), .A3(n3588), .A4(n3587), .ZN(n3611)
         );
  AOI22_X1 U3674 ( .A1(n3592), .A2(\xmem_inst/mem[41][1] ), .B1(n3591), .B2(
        \xmem_inst/mem[8][1] ), .ZN(n3596) );
  AOI22_X1 U3675 ( .A1(n3594), .A2(\xmem_inst/mem[19][1] ), .B1(n3593), .B2(
        \xmem_inst/mem[40][1] ), .ZN(n3595) );
  NAND2_X1 U3676 ( .A1(n3596), .A2(n3595), .ZN(n3610) );
  AOI22_X1 U3677 ( .A1(n3598), .A2(\xmem_inst/mem[0][1] ), .B1(n3597), .B2(
        \xmem_inst/mem[35][1] ), .ZN(n3608) );
  AOI22_X1 U3678 ( .A1(n3600), .A2(\xmem_inst/mem[21][1] ), .B1(n3599), .B2(
        \xmem_inst/mem[33][1] ), .ZN(n3607) );
  AOI22_X1 U3679 ( .A1(n3602), .A2(\xmem_inst/mem[32][1] ), .B1(n3601), .B2(
        \xmem_inst/mem[26][1] ), .ZN(n3606) );
  AOI22_X1 U3680 ( .A1(n3604), .A2(\xmem_inst/mem[4][1] ), .B1(n3603), .B2(
        \xmem_inst/mem[10][1] ), .ZN(n3605) );
  NAND4_X1 U3681 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(n3609)
         );
  NOR4_X1 U3682 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3639)
         );
  AOI22_X1 U3683 ( .A1(n3614), .A2(\xmem_inst/mem[23][1] ), .B1(n3613), .B2(
        \xmem_inst/mem[37][1] ), .ZN(n3638) );
  AOI22_X1 U3684 ( .A1(n3616), .A2(\xmem_inst/mem[14][1] ), .B1(n3615), .B2(
        \xmem_inst/mem[2][1] ), .ZN(n3623) );
  NAND2_X1 U3685 ( .A1(n3617), .A2(\xmem_inst/mem[42][1] ), .ZN(n3622) );
  NAND2_X1 U3686 ( .A1(n3618), .A2(\xmem_inst/mem[15][1] ), .ZN(n3621) );
  NAND2_X1 U3687 ( .A1(n3619), .A2(\xmem_inst/mem[9][1] ), .ZN(n3620) );
  AND4_X1 U3688 ( .A1(n3623), .A2(n3622), .A3(n3621), .A4(n3620), .ZN(n3637)
         );
  AOI22_X1 U3689 ( .A1(n3625), .A2(\xmem_inst/mem[6][1] ), .B1(n3624), .B2(
        \xmem_inst/mem[11][1] ), .ZN(n3635) );
  AOI22_X1 U3690 ( .A1(n3627), .A2(\xmem_inst/mem[39][1] ), .B1(n3626), .B2(
        \xmem_inst/mem[3][1] ), .ZN(n3634) );
  AOI22_X1 U3691 ( .A1(n3629), .A2(\xmem_inst/mem[31][1] ), .B1(n3628), .B2(
        \xmem_inst/mem[1][1] ), .ZN(n3633) );
  AOI22_X1 U3692 ( .A1(n3631), .A2(\xmem_inst/mem[34][1] ), .B1(n3630), .B2(
        \xmem_inst/mem[30][1] ), .ZN(n3632) );
  AND4_X1 U3693 ( .A1(n3635), .A2(n3634), .A3(n3633), .A4(n3632), .ZN(n3636)
         );
  NAND4_X1 U3694 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n3636), .ZN(
        \xmem_inst/N278 ) );
  NAND2_X1 U3695 ( .A1(n3641), .A2(n294), .ZN(n3642) );
  XOR2_X1 U3696 ( .A(n3643), .B(n3642), .Z(n3644) );
  NAND2_X1 U3697 ( .A1(n3646), .A2(n3645), .ZN(n3647) );
  XNOR2_X1 U3698 ( .A(n3648), .B(n3647), .ZN(n3649) );
  INV_X1 U3699 ( .A(n3650), .ZN(n3655) );
  INV_X1 U3700 ( .A(n3651), .ZN(n3653) );
  NAND2_X1 U3701 ( .A1(n3653), .A2(n3652), .ZN(n3654) );
  XOR2_X1 U3702 ( .A(n3655), .B(n3654), .Z(n3656) );
  NAND2_X1 U3703 ( .A1(n302), .A2(n3671), .ZN(n3662) );
  NAND2_X1 U3704 ( .A1(n3662), .A2(n3670), .ZN(n3666) );
  NAND2_X1 U3705 ( .A1(n3664), .A2(n3663), .ZN(n3665) );
  XNOR2_X1 U3706 ( .A(n3666), .B(n3665), .ZN(n3667) );
  NAND2_X1 U3707 ( .A1(n3671), .A2(n3670), .ZN(n3672) );
  XOR2_X1 U3708 ( .A(n3673), .B(n3672), .Z(n3674) );
  NAND2_X1 U3709 ( .A1(n3657), .A2(n3674), .ZN(n3675) );
  OAI211_X1 U3710 ( .C1(n2223), .C2(n4139), .A(n3675), .B(n3681), .ZN(
        \mac_unit_inst/n136 ) );
  NAND2_X1 U3711 ( .A1(n236), .A2(n3676), .ZN(n3677) );
  XNOR2_X1 U3712 ( .A(n3678), .B(n3677), .ZN(n3679) );
  NAND3_X1 U3713 ( .A1(n3684), .A2(n3683), .A3(n3682), .ZN(\fmem_inst/N76 ) );
  NAND3_X1 U3714 ( .A1(n3686), .A2(n4012), .A3(n3685), .ZN(\fmem_inst/N71 ) );
  NAND3_X1 U3715 ( .A1(n3688), .A2(n3687), .A3(n3695), .ZN(\fmem_inst/N68 ) );
  AOI22_X1 U3716 ( .A1(n3690), .A2(n4074), .B1(n3689), .B2(fmem_addr[1]), .ZN(
        n3692) );
  NAND2_X1 U3717 ( .A1(n3691), .A2(n4069), .ZN(n3694) );
  NAND3_X1 U3718 ( .A1(n3692), .A2(n4012), .A3(n3694), .ZN(\fmem_inst/N67 ) );
  INV_X1 U3719 ( .A(n3693), .ZN(n3696) );
  NAND3_X1 U3720 ( .A1(n3696), .A2(n3695), .A3(n3694), .ZN(\fmem_inst/N66 ) );
  NAND2_X1 U3721 ( .A1(n3710), .A2(n4105), .ZN(n3897) );
  NOR2_X2 U3722 ( .A1(n3897), .A2(n3723), .ZN(n3698) );
  INV_X2 U3723 ( .A(n3699), .ZN(n3700) );
  OAI22_X1 U3724 ( .A1(n3700), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[0][0] ), 
        .B2(n3699), .ZN(n4145) );
  OAI22_X1 U3725 ( .A1(n3700), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[0][1] ), 
        .B2(n3698), .ZN(n4146) );
  OAI22_X1 U3726 ( .A1(n3700), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[0][2] ), 
        .B2(n3698), .ZN(n4147) );
  OAI22_X1 U3727 ( .A1(n3700), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[0][3] ), 
        .B2(n3698), .ZN(n4148) );
  OAI22_X1 U3728 ( .A1(n3700), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[0][4] ), 
        .B2(n3698), .ZN(n4149) );
  OAI22_X1 U3729 ( .A1(n3700), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[0][5] ), 
        .B2(n3698), .ZN(n4150) );
  OAI22_X1 U3730 ( .A1(n3700), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[0][6] ), 
        .B2(n3698), .ZN(n4151) );
  OAI22_X1 U3731 ( .A1(n3700), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[0][7] ), 
        .B2(n3698), .ZN(n4152) );
  OAI22_X1 U3732 ( .A1(n3700), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[0][8] ), 
        .B2(n3698), .ZN(n4153) );
  OAI22_X1 U3733 ( .A1(n3700), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[0][9] ), 
        .B2(n3698), .ZN(n4154) );
  OAI22_X1 U3734 ( .A1(n3700), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[0][10] ), .B2(n3698), .ZN(n4155) );
  OAI22_X1 U3735 ( .A1(n3700), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[0][11] ), .B2(n3698), .ZN(n4156) );
  OAI22_X1 U3736 ( .A1(n3700), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[0][12] ), .B2(n3698), .ZN(n4157) );
  OAI22_X1 U3737 ( .A1(n3700), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[0][13] ), .B2(n3698), .ZN(n4158) );
  OAI22_X1 U3738 ( .A1(n3700), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[0][14] ), .B2(n3698), .ZN(n4159) );
  OAI22_X1 U3739 ( .A1(n3700), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[0][15] ), .B2(n3699), .ZN(n4160) );
  OAI22_X1 U3740 ( .A1(n3700), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[0][16] ), .B2(n3698), .ZN(n4161) );
  OAI22_X1 U3741 ( .A1(n3700), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[0][17] ), .B2(n3698), .ZN(n4162) );
  OAI22_X1 U3742 ( .A1(n3700), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[0][18] ), .B2(n3698), .ZN(n4163) );
  OAI22_X1 U3743 ( .A1(n3700), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[0][19] ), .B2(n3699), .ZN(n4164) );
  OAI22_X1 U3744 ( .A1(n3700), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[0][20] ), .B2(n3698), .ZN(n4165) );
  OAI22_X1 U3745 ( .A1(n3700), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[0][21] ), .B2(n3698), .ZN(n4166) );
  OAI22_X1 U3746 ( .A1(n3700), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[0][22] ), .B2(n3699), .ZN(n4167) );
  OAI22_X1 U3747 ( .A1(n3700), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[0][23] ), .B2(n3699), .ZN(n4168) );
  OAI22_X1 U3748 ( .A1(n3700), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[0][24] ), .B2(n3699), .ZN(n4169) );
  OAI22_X1 U3749 ( .A1(n3700), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[0][25] ), .B2(n3698), .ZN(n4170) );
  OAI22_X1 U3750 ( .A1(n3700), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[0][26] ), .B2(n3699), .ZN(n4171) );
  OAI22_X1 U3751 ( .A1(n3700), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[0][27] ), .B2(n3698), .ZN(n4172) );
  OAI22_X1 U3752 ( .A1(n3700), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[0][28] ), .B2(n3699), .ZN(n4173) );
  OAI22_X1 U3753 ( .A1(n3700), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[0][29] ), .B2(n3698), .ZN(n4174) );
  OAI22_X1 U3754 ( .A1(n3700), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[0][30] ), .B2(n3699), .ZN(n4175) );
  OAI22_X1 U3755 ( .A1(n3700), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[0][31] ), .B2(n3699), .ZN(n4176) );
  NAND2_X1 U3756 ( .A1(n3714), .A2(n4105), .ZN(n3933) );
  NOR2_X2 U3757 ( .A1(n3933), .A2(n3723), .ZN(n3701) );
  INV_X2 U3758 ( .A(n3702), .ZN(n3703) );
  OAI22_X1 U3759 ( .A1(n3703), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[1][0] ), 
        .B2(n3702), .ZN(n4177) );
  OAI22_X1 U3760 ( .A1(n3703), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[1][1] ), 
        .B2(n3701), .ZN(n4178) );
  OAI22_X1 U3761 ( .A1(n3703), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[1][2] ), 
        .B2(n3701), .ZN(n4179) );
  OAI22_X1 U3762 ( .A1(n3703), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[1][3] ), 
        .B2(n3701), .ZN(n4180) );
  OAI22_X1 U3763 ( .A1(n3703), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[1][4] ), 
        .B2(n3701), .ZN(n4181) );
  OAI22_X1 U3764 ( .A1(n3703), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[1][5] ), 
        .B2(n3701), .ZN(n4182) );
  OAI22_X1 U3765 ( .A1(n3703), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[1][6] ), 
        .B2(n3701), .ZN(n4183) );
  OAI22_X1 U3766 ( .A1(n3703), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[1][7] ), 
        .B2(n3701), .ZN(n4184) );
  OAI22_X1 U3767 ( .A1(n3703), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[1][8] ), 
        .B2(n3701), .ZN(n4185) );
  OAI22_X1 U3768 ( .A1(n3703), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[1][9] ), 
        .B2(n3701), .ZN(n4186) );
  OAI22_X1 U3769 ( .A1(n3703), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[1][10] ), .B2(n3701), .ZN(n4187) );
  OAI22_X1 U3770 ( .A1(n3703), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[1][11] ), .B2(n3701), .ZN(n4188) );
  OAI22_X1 U3771 ( .A1(n3703), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[1][12] ), .B2(n3701), .ZN(n4189) );
  OAI22_X1 U3772 ( .A1(n3703), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[1][13] ), .B2(n3701), .ZN(n4190) );
  OAI22_X1 U3773 ( .A1(n3703), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[1][14] ), .B2(n3701), .ZN(n4191) );
  OAI22_X1 U3774 ( .A1(n3703), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[1][15] ), .B2(n3702), .ZN(n4192) );
  OAI22_X1 U3775 ( .A1(n3703), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[1][16] ), .B2(n3701), .ZN(n4193) );
  OAI22_X1 U3776 ( .A1(n3703), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[1][17] ), .B2(n3701), .ZN(n4194) );
  OAI22_X1 U3777 ( .A1(n3703), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[1][18] ), .B2(n3701), .ZN(n4195) );
  OAI22_X1 U3778 ( .A1(n3703), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[1][19] ), .B2(n3702), .ZN(n4196) );
  OAI22_X1 U3779 ( .A1(n3703), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[1][20] ), .B2(n3701), .ZN(n4197) );
  OAI22_X1 U3780 ( .A1(n3703), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[1][21] ), .B2(n3701), .ZN(n4198) );
  OAI22_X1 U3781 ( .A1(n3703), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[1][22] ), .B2(n3702), .ZN(n4199) );
  OAI22_X1 U3782 ( .A1(n3703), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[1][23] ), .B2(n3702), .ZN(n4200) );
  OAI22_X1 U3783 ( .A1(n3703), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[1][24] ), .B2(n3702), .ZN(n4201) );
  OAI22_X1 U3784 ( .A1(n3703), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[1][25] ), .B2(n3701), .ZN(n4202) );
  OAI22_X1 U3785 ( .A1(n3703), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[1][26] ), .B2(n3702), .ZN(n4203) );
  OAI22_X1 U3786 ( .A1(n3703), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[1][27] ), .B2(n3701), .ZN(n4204) );
  OAI22_X1 U3787 ( .A1(n3703), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[1][28] ), .B2(n3702), .ZN(n4205) );
  OAI22_X1 U3788 ( .A1(n3703), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[1][29] ), .B2(n3701), .ZN(n4206) );
  OAI22_X1 U3789 ( .A1(n3703), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[1][30] ), .B2(n3702), .ZN(n4207) );
  OAI22_X1 U3790 ( .A1(n3703), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[1][31] ), .B2(n3702), .ZN(n4208) );
  NAND2_X1 U3791 ( .A1(n3718), .A2(n4105), .ZN(n3970) );
  NOR2_X2 U3792 ( .A1(n3970), .A2(n3723), .ZN(n3704) );
  INV_X2 U3793 ( .A(n3705), .ZN(n3706) );
  OAI22_X1 U3794 ( .A1(n3706), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[2][0] ), 
        .B2(n3705), .ZN(n4209) );
  OAI22_X1 U3795 ( .A1(n3706), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[2][1] ), 
        .B2(n3704), .ZN(n4210) );
  OAI22_X1 U3796 ( .A1(n3706), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[2][2] ), 
        .B2(n3704), .ZN(n4211) );
  OAI22_X1 U3797 ( .A1(n3706), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[2][3] ), 
        .B2(n3704), .ZN(n4212) );
  OAI22_X1 U3798 ( .A1(n3706), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[2][4] ), 
        .B2(n3704), .ZN(n4213) );
  OAI22_X1 U3799 ( .A1(n3706), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[2][5] ), 
        .B2(n3704), .ZN(n4214) );
  OAI22_X1 U3800 ( .A1(n3706), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[2][6] ), 
        .B2(n3704), .ZN(n4215) );
  OAI22_X1 U3801 ( .A1(n3706), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[2][7] ), 
        .B2(n3704), .ZN(n4216) );
  OAI22_X1 U3802 ( .A1(n3706), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[2][8] ), 
        .B2(n3704), .ZN(n4217) );
  OAI22_X1 U3803 ( .A1(n3706), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[2][9] ), 
        .B2(n3704), .ZN(n4218) );
  OAI22_X1 U3804 ( .A1(n3706), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[2][10] ), .B2(n3704), .ZN(n4219) );
  OAI22_X1 U3805 ( .A1(n3706), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[2][11] ), .B2(n3704), .ZN(n4220) );
  OAI22_X1 U3806 ( .A1(n3706), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[2][12] ), .B2(n3704), .ZN(n4221) );
  OAI22_X1 U3807 ( .A1(n3706), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[2][13] ), .B2(n3704), .ZN(n4222) );
  OAI22_X1 U3808 ( .A1(n3706), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[2][14] ), .B2(n3704), .ZN(n4223) );
  OAI22_X1 U3809 ( .A1(n3706), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[2][15] ), .B2(n3705), .ZN(n4224) );
  OAI22_X1 U3810 ( .A1(n3706), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[2][16] ), .B2(n3704), .ZN(n4225) );
  OAI22_X1 U3811 ( .A1(n3706), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[2][17] ), .B2(n3704), .ZN(n4226) );
  OAI22_X1 U3812 ( .A1(n3706), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[2][18] ), .B2(n3704), .ZN(n4227) );
  OAI22_X1 U3813 ( .A1(n3706), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[2][19] ), .B2(n3705), .ZN(n4228) );
  OAI22_X1 U3814 ( .A1(n3706), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[2][20] ), .B2(n3704), .ZN(n4229) );
  OAI22_X1 U3815 ( .A1(n3706), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[2][21] ), .B2(n3704), .ZN(n4230) );
  OAI22_X1 U3816 ( .A1(n3706), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[2][22] ), .B2(n3705), .ZN(n4231) );
  OAI22_X1 U3817 ( .A1(n3706), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[2][23] ), .B2(n3705), .ZN(n4232) );
  OAI22_X1 U3818 ( .A1(n3706), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[2][24] ), .B2(n3705), .ZN(n4233) );
  OAI22_X1 U3819 ( .A1(n3706), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[2][25] ), .B2(n3704), .ZN(n4234) );
  OAI22_X1 U3820 ( .A1(n3706), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[2][26] ), .B2(n3705), .ZN(n4235) );
  OAI22_X1 U3821 ( .A1(n3706), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[2][27] ), .B2(n3704), .ZN(n4236) );
  OAI22_X1 U3822 ( .A1(n3706), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[2][28] ), .B2(n3705), .ZN(n4237) );
  OAI22_X1 U3823 ( .A1(n3706), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[2][29] ), .B2(n3704), .ZN(n4238) );
  OAI22_X1 U3824 ( .A1(n3706), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[2][30] ), .B2(n3705), .ZN(n4239) );
  OAI22_X1 U3825 ( .A1(n3706), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[2][31] ), .B2(n3705), .ZN(n4240) );
  NAND2_X1 U3826 ( .A1(n3722), .A2(n4105), .ZN(n3873) );
  NOR2_X2 U3827 ( .A1(n3873), .A2(n3723), .ZN(n3707) );
  INV_X2 U3828 ( .A(n3708), .ZN(n3709) );
  OAI22_X1 U3829 ( .A1(n3709), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[3][0] ), 
        .B2(n3708), .ZN(n4241) );
  OAI22_X1 U3830 ( .A1(n3709), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[3][1] ), 
        .B2(n3707), .ZN(n4242) );
  OAI22_X1 U3831 ( .A1(n3709), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[3][2] ), 
        .B2(n3707), .ZN(n4243) );
  OAI22_X1 U3832 ( .A1(n3709), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[3][3] ), 
        .B2(n3707), .ZN(n4244) );
  OAI22_X1 U3833 ( .A1(n3709), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[3][4] ), 
        .B2(n3707), .ZN(n4245) );
  OAI22_X1 U3834 ( .A1(n3709), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[3][5] ), 
        .B2(n3707), .ZN(n4246) );
  OAI22_X1 U3835 ( .A1(n3709), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[3][6] ), 
        .B2(n3707), .ZN(n4247) );
  OAI22_X1 U3836 ( .A1(n3709), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[3][7] ), 
        .B2(n3707), .ZN(n4248) );
  OAI22_X1 U3837 ( .A1(n3709), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[3][8] ), 
        .B2(n3707), .ZN(n4249) );
  OAI22_X1 U3838 ( .A1(n3709), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[3][9] ), 
        .B2(n3707), .ZN(n4250) );
  OAI22_X1 U3839 ( .A1(n3709), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[3][10] ), .B2(n3707), .ZN(n4251) );
  OAI22_X1 U3840 ( .A1(n3709), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[3][11] ), .B2(n3707), .ZN(n4252) );
  OAI22_X1 U3841 ( .A1(n3709), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[3][12] ), .B2(n3707), .ZN(n4253) );
  OAI22_X1 U3842 ( .A1(n3709), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[3][13] ), .B2(n3707), .ZN(n4254) );
  OAI22_X1 U3843 ( .A1(n3709), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[3][14] ), .B2(n3707), .ZN(n4255) );
  OAI22_X1 U3844 ( .A1(n3709), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[3][15] ), .B2(n3708), .ZN(n4256) );
  OAI22_X1 U3845 ( .A1(n3709), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[3][16] ), .B2(n3707), .ZN(n4257) );
  OAI22_X1 U3846 ( .A1(n3709), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[3][17] ), .B2(n3707), .ZN(n4258) );
  OAI22_X1 U3847 ( .A1(n3709), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[3][18] ), .B2(n3707), .ZN(n4259) );
  OAI22_X1 U3848 ( .A1(n3709), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[3][19] ), .B2(n3708), .ZN(n4260) );
  OAI22_X1 U3849 ( .A1(n3709), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[3][20] ), .B2(n3707), .ZN(n4261) );
  OAI22_X1 U3850 ( .A1(n3709), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[3][21] ), .B2(n3707), .ZN(n4262) );
  OAI22_X1 U3851 ( .A1(n3709), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[3][22] ), .B2(n3708), .ZN(n4263) );
  OAI22_X1 U3852 ( .A1(n3709), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[3][23] ), .B2(n3708), .ZN(n4264) );
  OAI22_X1 U3853 ( .A1(n3709), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[3][24] ), .B2(n3708), .ZN(n4265) );
  OAI22_X1 U3854 ( .A1(n3709), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[3][25] ), .B2(n3707), .ZN(n4266) );
  OAI22_X1 U3855 ( .A1(n3709), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[3][26] ), .B2(n3708), .ZN(n4267) );
  OAI22_X1 U3856 ( .A1(n3709), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[3][27] ), .B2(n3707), .ZN(n4268) );
  OAI22_X1 U3857 ( .A1(n3709), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[3][28] ), .B2(n3708), .ZN(n4269) );
  OAI22_X1 U3858 ( .A1(n3709), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[3][29] ), .B2(n3707), .ZN(n4270) );
  OAI22_X1 U3859 ( .A1(n3709), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[3][30] ), .B2(n3708), .ZN(n4271) );
  OAI22_X1 U3860 ( .A1(n3709), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[3][31] ), .B2(n3708), .ZN(n4272) );
  NAND2_X1 U3861 ( .A1(xmem_addr[2]), .A2(n3710), .ZN(n3878) );
  NOR2_X2 U3862 ( .A1(n3878), .A2(n3723), .ZN(n3711) );
  INV_X2 U3863 ( .A(n3712), .ZN(n3713) );
  OAI22_X1 U3864 ( .A1(n3713), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[4][0] ), 
        .B2(n3712), .ZN(n4273) );
  OAI22_X1 U3865 ( .A1(n3713), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[4][1] ), 
        .B2(n3711), .ZN(n4274) );
  OAI22_X1 U3866 ( .A1(n3713), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[4][2] ), 
        .B2(n3711), .ZN(n4275) );
  OAI22_X1 U3867 ( .A1(n3713), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[4][3] ), 
        .B2(n3711), .ZN(n4276) );
  OAI22_X1 U3868 ( .A1(n3713), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[4][4] ), 
        .B2(n3711), .ZN(n4277) );
  OAI22_X1 U3869 ( .A1(n3713), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[4][5] ), 
        .B2(n3711), .ZN(n4278) );
  OAI22_X1 U3870 ( .A1(n3713), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[4][6] ), 
        .B2(n3711), .ZN(n4279) );
  OAI22_X1 U3871 ( .A1(n3713), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[4][7] ), 
        .B2(n3711), .ZN(n4280) );
  OAI22_X1 U3872 ( .A1(n3713), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[4][8] ), 
        .B2(n3711), .ZN(n4281) );
  OAI22_X1 U3873 ( .A1(n3713), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[4][9] ), 
        .B2(n3711), .ZN(n4282) );
  OAI22_X1 U3874 ( .A1(n3713), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[4][10] ), .B2(n3711), .ZN(n4283) );
  OAI22_X1 U3875 ( .A1(n3713), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[4][11] ), .B2(n3711), .ZN(n4284) );
  OAI22_X1 U3876 ( .A1(n3713), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[4][12] ), .B2(n3711), .ZN(n4285) );
  OAI22_X1 U3877 ( .A1(n3713), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[4][13] ), .B2(n3711), .ZN(n4286) );
  OAI22_X1 U3878 ( .A1(n3713), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[4][14] ), .B2(n3711), .ZN(n4287) );
  OAI22_X1 U3879 ( .A1(n3713), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[4][15] ), .B2(n3712), .ZN(n4288) );
  OAI22_X1 U3880 ( .A1(n3713), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[4][16] ), .B2(n3711), .ZN(n4289) );
  OAI22_X1 U3881 ( .A1(n3713), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[4][17] ), .B2(n3711), .ZN(n4290) );
  OAI22_X1 U3882 ( .A1(n3713), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[4][18] ), .B2(n3711), .ZN(n4291) );
  OAI22_X1 U3883 ( .A1(n3713), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[4][19] ), .B2(n3712), .ZN(n4292) );
  OAI22_X1 U3884 ( .A1(n3713), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[4][20] ), .B2(n3711), .ZN(n4293) );
  OAI22_X1 U3885 ( .A1(n3713), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[4][21] ), .B2(n3711), .ZN(n4294) );
  OAI22_X1 U3886 ( .A1(n3713), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[4][22] ), .B2(n3712), .ZN(n4295) );
  OAI22_X1 U3887 ( .A1(n3713), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[4][23] ), .B2(n3712), .ZN(n4296) );
  OAI22_X1 U3888 ( .A1(n3713), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[4][24] ), .B2(n3712), .ZN(n4297) );
  OAI22_X1 U3889 ( .A1(n3713), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[4][25] ), .B2(n3711), .ZN(n4298) );
  OAI22_X1 U3890 ( .A1(n3713), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[4][26] ), .B2(n3712), .ZN(n4299) );
  OAI22_X1 U3891 ( .A1(n3713), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[4][27] ), .B2(n3711), .ZN(n4300) );
  OAI22_X1 U3892 ( .A1(n3713), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[4][28] ), .B2(n3712), .ZN(n4301) );
  OAI22_X1 U3893 ( .A1(n3713), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[4][29] ), .B2(n3711), .ZN(n4302) );
  OAI22_X1 U3894 ( .A1(n3713), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[4][30] ), .B2(n3712), .ZN(n4303) );
  OAI22_X1 U3895 ( .A1(n3713), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[4][31] ), .B2(n3712), .ZN(n4304) );
  NAND2_X1 U3896 ( .A1(xmem_addr[2]), .A2(n3714), .ZN(n3882) );
  NOR2_X2 U3897 ( .A1(n3882), .A2(n3723), .ZN(n3715) );
  INV_X2 U3898 ( .A(n3716), .ZN(n3717) );
  OAI22_X1 U3899 ( .A1(n3717), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[5][0] ), 
        .B2(n3716), .ZN(n4305) );
  OAI22_X1 U3900 ( .A1(n3717), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[5][1] ), 
        .B2(n3715), .ZN(n4306) );
  OAI22_X1 U3901 ( .A1(n3717), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[5][2] ), 
        .B2(n3715), .ZN(n4307) );
  OAI22_X1 U3902 ( .A1(n3717), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[5][3] ), 
        .B2(n3715), .ZN(n4308) );
  OAI22_X1 U3903 ( .A1(n3717), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[5][4] ), 
        .B2(n3715), .ZN(n4309) );
  OAI22_X1 U3904 ( .A1(n3717), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[5][5] ), 
        .B2(n3715), .ZN(n4310) );
  OAI22_X1 U3905 ( .A1(n3717), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[5][6] ), 
        .B2(n3715), .ZN(n4311) );
  OAI22_X1 U3906 ( .A1(n3717), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[5][7] ), 
        .B2(n3715), .ZN(n4312) );
  OAI22_X1 U3907 ( .A1(n3717), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[5][8] ), 
        .B2(n3715), .ZN(n4313) );
  OAI22_X1 U3908 ( .A1(n3717), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[5][9] ), 
        .B2(n3715), .ZN(n4314) );
  OAI22_X1 U3909 ( .A1(n3717), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[5][10] ), .B2(n3715), .ZN(n4315) );
  OAI22_X1 U3910 ( .A1(n3717), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[5][11] ), .B2(n3715), .ZN(n4316) );
  OAI22_X1 U3911 ( .A1(n3717), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[5][12] ), .B2(n3715), .ZN(n4317) );
  OAI22_X1 U3912 ( .A1(n3717), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[5][13] ), .B2(n3715), .ZN(n4318) );
  OAI22_X1 U3913 ( .A1(n3717), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[5][14] ), .B2(n3715), .ZN(n4319) );
  OAI22_X1 U3914 ( .A1(n3717), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[5][15] ), .B2(n3716), .ZN(n4320) );
  OAI22_X1 U3915 ( .A1(n3717), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[5][16] ), .B2(n3715), .ZN(n4321) );
  OAI22_X1 U3916 ( .A1(n3717), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[5][17] ), .B2(n3715), .ZN(n4322) );
  OAI22_X1 U3917 ( .A1(n3717), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[5][18] ), .B2(n3715), .ZN(n4323) );
  OAI22_X1 U3918 ( .A1(n3717), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[5][19] ), .B2(n3716), .ZN(n4324) );
  OAI22_X1 U3919 ( .A1(n3717), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[5][20] ), .B2(n3715), .ZN(n4325) );
  OAI22_X1 U3920 ( .A1(n3717), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[5][21] ), .B2(n3715), .ZN(n4326) );
  OAI22_X1 U3921 ( .A1(n3717), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[5][22] ), .B2(n3716), .ZN(n4327) );
  OAI22_X1 U3922 ( .A1(n3717), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[5][23] ), .B2(n3716), .ZN(n4328) );
  OAI22_X1 U3923 ( .A1(n3717), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[5][24] ), .B2(n3716), .ZN(n4329) );
  OAI22_X1 U3924 ( .A1(n3717), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[5][25] ), .B2(n3715), .ZN(n4330) );
  OAI22_X1 U3925 ( .A1(n3717), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[5][26] ), .B2(n3716), .ZN(n4331) );
  OAI22_X1 U3926 ( .A1(n3717), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[5][27] ), .B2(n3715), .ZN(n4332) );
  OAI22_X1 U3927 ( .A1(n3717), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[5][28] ), .B2(n3716), .ZN(n4333) );
  OAI22_X1 U3928 ( .A1(n3717), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[5][29] ), .B2(n3715), .ZN(n4334) );
  OAI22_X1 U3929 ( .A1(n3717), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[5][30] ), .B2(n3716), .ZN(n4335) );
  OAI22_X1 U3930 ( .A1(n3717), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[5][31] ), .B2(n3716), .ZN(n4336) );
  NAND2_X1 U3931 ( .A1(xmem_addr[2]), .A2(n3718), .ZN(n3886) );
  NOR2_X2 U3932 ( .A1(n3886), .A2(n3723), .ZN(n3719) );
  INV_X2 U3933 ( .A(n3720), .ZN(n3721) );
  OAI22_X1 U3934 ( .A1(n3721), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[6][0] ), 
        .B2(n3720), .ZN(n4337) );
  OAI22_X1 U3935 ( .A1(n3721), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[6][1] ), 
        .B2(n3719), .ZN(n4338) );
  OAI22_X1 U3936 ( .A1(n3721), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[6][2] ), 
        .B2(n3719), .ZN(n4339) );
  OAI22_X1 U3937 ( .A1(n3721), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[6][3] ), 
        .B2(n3719), .ZN(n4340) );
  OAI22_X1 U3938 ( .A1(n3721), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[6][4] ), 
        .B2(n3719), .ZN(n4341) );
  OAI22_X1 U3939 ( .A1(n3721), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[6][5] ), 
        .B2(n3719), .ZN(n4342) );
  OAI22_X1 U3940 ( .A1(n3721), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[6][6] ), 
        .B2(n3719), .ZN(n4343) );
  OAI22_X1 U3941 ( .A1(n3721), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[6][7] ), 
        .B2(n3719), .ZN(n4344) );
  OAI22_X1 U3942 ( .A1(n3721), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[6][8] ), 
        .B2(n3719), .ZN(n4345) );
  OAI22_X1 U3943 ( .A1(n3721), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[6][9] ), 
        .B2(n3719), .ZN(n4346) );
  OAI22_X1 U3944 ( .A1(n3721), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[6][10] ), .B2(n3719), .ZN(n4347) );
  OAI22_X1 U3945 ( .A1(n3721), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[6][11] ), .B2(n3719), .ZN(n4348) );
  OAI22_X1 U3946 ( .A1(n3721), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[6][12] ), .B2(n3719), .ZN(n4349) );
  OAI22_X1 U3947 ( .A1(n3721), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[6][13] ), .B2(n3719), .ZN(n4350) );
  OAI22_X1 U3948 ( .A1(n3721), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[6][14] ), .B2(n3719), .ZN(n4351) );
  OAI22_X1 U3949 ( .A1(n3721), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[6][15] ), .B2(n3720), .ZN(n4352) );
  OAI22_X1 U3950 ( .A1(n3721), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[6][16] ), .B2(n3719), .ZN(n4353) );
  OAI22_X1 U3951 ( .A1(n3721), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[6][17] ), .B2(n3719), .ZN(n4354) );
  OAI22_X1 U3952 ( .A1(n3721), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[6][18] ), .B2(n3719), .ZN(n4355) );
  OAI22_X1 U3953 ( .A1(n3721), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[6][19] ), .B2(n3720), .ZN(n4356) );
  OAI22_X1 U3954 ( .A1(n3721), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[6][20] ), .B2(n3719), .ZN(n4357) );
  OAI22_X1 U3955 ( .A1(n3721), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[6][21] ), .B2(n3719), .ZN(n4358) );
  OAI22_X1 U3956 ( .A1(n3721), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[6][22] ), .B2(n3720), .ZN(n4359) );
  OAI22_X1 U3957 ( .A1(n3721), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[6][23] ), .B2(n3720), .ZN(n4360) );
  OAI22_X1 U3958 ( .A1(n3721), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[6][24] ), .B2(n3720), .ZN(n4361) );
  OAI22_X1 U3959 ( .A1(n3721), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[6][25] ), .B2(n3719), .ZN(n4362) );
  OAI22_X1 U3960 ( .A1(n3721), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[6][26] ), .B2(n3720), .ZN(n4363) );
  OAI22_X1 U3961 ( .A1(n3721), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[6][27] ), .B2(n3719), .ZN(n4364) );
  OAI22_X1 U3962 ( .A1(n3721), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[6][28] ), .B2(n3720), .ZN(n4365) );
  OAI22_X1 U3963 ( .A1(n3721), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[6][29] ), .B2(n3719), .ZN(n4366) );
  OAI22_X1 U3964 ( .A1(n3721), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[6][30] ), .B2(n3720), .ZN(n4367) );
  OAI22_X1 U3965 ( .A1(n3721), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[6][31] ), .B2(n3720), .ZN(n4368) );
  NAND2_X1 U3966 ( .A1(n3722), .A2(xmem_addr[2]), .ZN(n3891) );
  NOR2_X2 U3967 ( .A1(n3891), .A2(n3723), .ZN(n3725) );
  INV_X2 U3968 ( .A(n3726), .ZN(n3727) );
  OAI22_X1 U3969 ( .A1(n3727), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[7][0] ), 
        .B2(n3725), .ZN(n4369) );
  OAI22_X1 U3970 ( .A1(n3727), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[7][1] ), 
        .B2(n3725), .ZN(n4370) );
  OAI22_X1 U3971 ( .A1(n3727), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[7][2] ), 
        .B2(n3725), .ZN(n4371) );
  OAI22_X1 U3972 ( .A1(n3727), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[7][3] ), 
        .B2(n3725), .ZN(n4372) );
  OAI22_X1 U3973 ( .A1(n3727), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[7][4] ), 
        .B2(n3725), .ZN(n4373) );
  OAI22_X1 U3974 ( .A1(n3727), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[7][5] ), 
        .B2(n3725), .ZN(n4374) );
  OAI22_X1 U3975 ( .A1(n3727), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[7][6] ), 
        .B2(n3725), .ZN(n4375) );
  OAI22_X1 U3976 ( .A1(n3727), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[7][7] ), 
        .B2(n3725), .ZN(n4376) );
  OAI22_X1 U3977 ( .A1(n3727), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[7][8] ), 
        .B2(n3725), .ZN(n4377) );
  OAI22_X1 U3978 ( .A1(n3727), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[7][9] ), 
        .B2(n3725), .ZN(n4378) );
  OAI22_X1 U3979 ( .A1(n3727), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[7][10] ), .B2(n3725), .ZN(n4379) );
  OAI22_X1 U3980 ( .A1(n3727), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[7][11] ), .B2(n3725), .ZN(n4380) );
  OAI22_X1 U3981 ( .A1(n3727), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[7][12] ), .B2(n3725), .ZN(n4381) );
  OAI22_X1 U3982 ( .A1(n3727), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[7][13] ), .B2(n3725), .ZN(n4382) );
  OAI22_X1 U3983 ( .A1(n3727), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[7][14] ), .B2(n3725), .ZN(n4383) );
  OAI22_X1 U3984 ( .A1(n3727), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[7][15] ), .B2(n3726), .ZN(n4384) );
  OAI22_X1 U3985 ( .A1(n3727), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[7][16] ), .B2(n3725), .ZN(n4385) );
  OAI22_X1 U3986 ( .A1(n3727), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[7][17] ), .B2(n3725), .ZN(n4386) );
  OAI22_X1 U3987 ( .A1(n3727), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[7][18] ), .B2(n3725), .ZN(n4387) );
  OAI22_X1 U3988 ( .A1(n3727), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[7][19] ), .B2(n3726), .ZN(n4388) );
  OAI22_X1 U3989 ( .A1(n3727), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[7][20] ), .B2(n3726), .ZN(n3724) );
  INV_X1 U3990 ( .A(n3724), .ZN(\xmem_inst/n2686 ) );
  OAI22_X1 U3991 ( .A1(n3727), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[7][21] ), .B2(n3725), .ZN(n4389) );
  OAI22_X1 U3992 ( .A1(n3727), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[7][22] ), .B2(n3726), .ZN(n4390) );
  OAI22_X1 U3993 ( .A1(n3727), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[7][23] ), .B2(n3726), .ZN(n4391) );
  OAI22_X1 U3994 ( .A1(n3727), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[7][24] ), .B2(n3726), .ZN(n4392) );
  OAI22_X1 U3995 ( .A1(n3727), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[7][25] ), .B2(n3725), .ZN(n4393) );
  OAI22_X1 U3996 ( .A1(n3727), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[7][26] ), .B2(n3726), .ZN(n4394) );
  OAI22_X1 U3997 ( .A1(n3727), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[7][27] ), .B2(n3725), .ZN(n4395) );
  OAI22_X1 U3998 ( .A1(n3727), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[7][28] ), .B2(n3726), .ZN(n4396) );
  OAI22_X1 U3999 ( .A1(n3727), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[7][29] ), .B2(n3725), .ZN(n4397) );
  OAI22_X1 U4000 ( .A1(n3727), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[7][30] ), .B2(n3726), .ZN(n4398) );
  OAI22_X1 U4001 ( .A1(n3727), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[7][31] ), .B2(n3726), .ZN(n4399) );
  NOR2_X2 U4002 ( .A1(n3897), .A2(n3750), .ZN(n3729) );
  INV_X2 U4003 ( .A(n3730), .ZN(n3731) );
  OAI22_X1 U4004 ( .A1(n3731), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[8][0] ), 
        .B2(n3730), .ZN(n4400) );
  OAI22_X1 U4005 ( .A1(n3731), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[8][1] ), 
        .B2(n3729), .ZN(n4401) );
  OAI22_X1 U4006 ( .A1(n3731), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[8][2] ), 
        .B2(n3729), .ZN(n4402) );
  OAI22_X1 U4007 ( .A1(n3731), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[8][3] ), 
        .B2(n3729), .ZN(n4403) );
  OAI22_X1 U4008 ( .A1(n3731), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[8][4] ), 
        .B2(n3729), .ZN(n4404) );
  OAI22_X1 U4009 ( .A1(n3731), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[8][5] ), 
        .B2(n3729), .ZN(n4405) );
  OAI22_X1 U4010 ( .A1(n3731), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[8][6] ), 
        .B2(n3729), .ZN(n4406) );
  OAI22_X1 U4011 ( .A1(n3731), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[8][7] ), 
        .B2(n3729), .ZN(n4407) );
  OAI22_X1 U4012 ( .A1(n3731), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[8][8] ), 
        .B2(n3729), .ZN(n4408) );
  OAI22_X1 U4013 ( .A1(n3731), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[8][9] ), 
        .B2(n3729), .ZN(n4409) );
  OAI22_X1 U4014 ( .A1(n3731), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[8][10] ), .B2(n3729), .ZN(n4410) );
  OAI22_X1 U4015 ( .A1(n3731), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[8][11] ), .B2(n3729), .ZN(n4411) );
  OAI22_X1 U4016 ( .A1(n3731), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[8][12] ), .B2(n3729), .ZN(n4412) );
  OAI22_X1 U4017 ( .A1(n3731), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[8][13] ), .B2(n3729), .ZN(n4413) );
  OAI22_X1 U4018 ( .A1(n3731), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[8][14] ), .B2(n3729), .ZN(n4414) );
  OAI22_X1 U4019 ( .A1(n3731), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[8][15] ), .B2(n3730), .ZN(n4415) );
  OAI22_X1 U4020 ( .A1(n3731), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[8][16] ), .B2(n3729), .ZN(n4416) );
  OAI22_X1 U4021 ( .A1(n3731), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[8][17] ), .B2(n3729), .ZN(n4417) );
  OAI22_X1 U4022 ( .A1(n3731), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[8][18] ), .B2(n3729), .ZN(n4418) );
  OAI22_X1 U4023 ( .A1(n3731), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[8][19] ), .B2(n3730), .ZN(n4419) );
  OAI22_X1 U4024 ( .A1(n3731), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[8][20] ), .B2(n3729), .ZN(n4420) );
  OAI22_X1 U4025 ( .A1(n3731), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[8][21] ), .B2(n3729), .ZN(n4421) );
  OAI22_X1 U4026 ( .A1(n3731), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[8][22] ), .B2(n3730), .ZN(n4422) );
  OAI22_X1 U4027 ( .A1(n3731), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[8][23] ), .B2(n3730), .ZN(n4423) );
  OAI22_X1 U4028 ( .A1(n3731), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[8][24] ), .B2(n3730), .ZN(n4424) );
  OAI22_X1 U4029 ( .A1(n3731), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[8][25] ), .B2(n3729), .ZN(n4425) );
  OAI22_X1 U4030 ( .A1(n3731), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[8][26] ), .B2(n3730), .ZN(n4426) );
  OAI22_X1 U4031 ( .A1(n3731), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[8][27] ), .B2(n3729), .ZN(n4427) );
  OAI22_X1 U4032 ( .A1(n3731), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[8][28] ), .B2(n3730), .ZN(n4428) );
  OAI22_X1 U4033 ( .A1(n3731), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[8][29] ), .B2(n3729), .ZN(n4429) );
  OAI22_X1 U4034 ( .A1(n3731), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[8][30] ), .B2(n3730), .ZN(n4430) );
  OAI22_X1 U4035 ( .A1(n3731), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[8][31] ), .B2(n3730), .ZN(n4431) );
  NOR2_X2 U4036 ( .A1(n3933), .A2(n3750), .ZN(n3732) );
  INV_X2 U4037 ( .A(n3733), .ZN(n3734) );
  OAI22_X1 U4038 ( .A1(n3734), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[9][0] ), 
        .B2(n3733), .ZN(n4432) );
  OAI22_X1 U4039 ( .A1(n3734), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[9][1] ), 
        .B2(n3732), .ZN(n4433) );
  OAI22_X1 U4040 ( .A1(n3734), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[9][2] ), 
        .B2(n3732), .ZN(n4434) );
  OAI22_X1 U4041 ( .A1(n3734), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[9][3] ), 
        .B2(n3732), .ZN(n4435) );
  OAI22_X1 U4042 ( .A1(n3734), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[9][4] ), 
        .B2(n3732), .ZN(n4436) );
  OAI22_X1 U4043 ( .A1(n3734), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[9][5] ), 
        .B2(n3732), .ZN(n4437) );
  OAI22_X1 U4044 ( .A1(n3734), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[9][6] ), 
        .B2(n3732), .ZN(n4438) );
  OAI22_X1 U4045 ( .A1(n3734), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[9][7] ), 
        .B2(n3732), .ZN(n4439) );
  OAI22_X1 U4046 ( .A1(n3734), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[9][8] ), 
        .B2(n3732), .ZN(n4440) );
  OAI22_X1 U4047 ( .A1(n3734), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[9][9] ), 
        .B2(n3732), .ZN(n4441) );
  OAI22_X1 U4048 ( .A1(n3734), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[9][10] ), .B2(n3732), .ZN(n4442) );
  OAI22_X1 U4049 ( .A1(n3734), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[9][11] ), .B2(n3732), .ZN(n4443) );
  OAI22_X1 U4050 ( .A1(n3734), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[9][12] ), .B2(n3732), .ZN(n4444) );
  OAI22_X1 U4051 ( .A1(n3734), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[9][13] ), .B2(n3732), .ZN(n4445) );
  OAI22_X1 U4052 ( .A1(n3734), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[9][14] ), .B2(n3732), .ZN(n4446) );
  OAI22_X1 U4053 ( .A1(n3734), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[9][15] ), .B2(n3733), .ZN(n4447) );
  OAI22_X1 U4054 ( .A1(n3734), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[9][16] ), .B2(n3732), .ZN(n4448) );
  OAI22_X1 U4055 ( .A1(n3734), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[9][17] ), .B2(n3732), .ZN(n4449) );
  OAI22_X1 U4056 ( .A1(n3734), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[9][18] ), .B2(n3732), .ZN(n4450) );
  OAI22_X1 U4057 ( .A1(n3734), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[9][19] ), .B2(n3733), .ZN(n4451) );
  OAI22_X1 U4058 ( .A1(n3734), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[9][20] ), .B2(n3732), .ZN(n4452) );
  OAI22_X1 U4059 ( .A1(n3734), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[9][21] ), .B2(n3732), .ZN(n4453) );
  OAI22_X1 U4060 ( .A1(n3734), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[9][22] ), .B2(n3733), .ZN(n4454) );
  OAI22_X1 U4061 ( .A1(n3734), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[9][23] ), .B2(n3733), .ZN(n4455) );
  OAI22_X1 U4062 ( .A1(n3734), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[9][24] ), .B2(n3733), .ZN(n4456) );
  OAI22_X1 U4063 ( .A1(n3734), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[9][25] ), .B2(n3732), .ZN(n4457) );
  OAI22_X1 U4064 ( .A1(n3734), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[9][26] ), .B2(n3733), .ZN(n4458) );
  OAI22_X1 U4065 ( .A1(n3734), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[9][27] ), .B2(n3732), .ZN(n4459) );
  OAI22_X1 U4066 ( .A1(n3734), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[9][28] ), .B2(n3733), .ZN(n4460) );
  OAI22_X1 U4067 ( .A1(n3734), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[9][29] ), .B2(n3732), .ZN(n4461) );
  OAI22_X1 U4068 ( .A1(n3734), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[9][30] ), .B2(n3733), .ZN(n4462) );
  OAI22_X1 U4069 ( .A1(n3734), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[9][31] ), .B2(n3733), .ZN(n4463) );
  NOR2_X2 U4070 ( .A1(n3970), .A2(n3750), .ZN(n3735) );
  INV_X2 U4071 ( .A(n3736), .ZN(n3737) );
  OAI22_X1 U4072 ( .A1(n3737), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[10][0] ), .B2(n3736), .ZN(n4464) );
  OAI22_X1 U4073 ( .A1(n3737), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[10][1] ), .B2(n3735), .ZN(n4465) );
  OAI22_X1 U4074 ( .A1(n3737), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[10][2] ), .B2(n3735), .ZN(n4466) );
  OAI22_X1 U4075 ( .A1(n3737), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[10][3] ), .B2(n3735), .ZN(n4467) );
  OAI22_X1 U4076 ( .A1(n3737), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[10][4] ), .B2(n3735), .ZN(n4468) );
  OAI22_X1 U4077 ( .A1(n3737), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[10][5] ), .B2(n3735), .ZN(n4469) );
  OAI22_X1 U4078 ( .A1(n3737), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[10][6] ), .B2(n3735), .ZN(n4470) );
  OAI22_X1 U4079 ( .A1(n3737), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[10][7] ), .B2(n3735), .ZN(n4471) );
  OAI22_X1 U4080 ( .A1(n3737), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[10][8] ), .B2(n3735), .ZN(n4472) );
  OAI22_X1 U4081 ( .A1(n3737), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[10][9] ), .B2(n3735), .ZN(n4473) );
  OAI22_X1 U4082 ( .A1(n3737), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[10][10] ), .B2(n3735), .ZN(n4474) );
  OAI22_X1 U4083 ( .A1(n3737), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[10][11] ), .B2(n3735), .ZN(n4475) );
  OAI22_X1 U4084 ( .A1(n3737), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[10][12] ), .B2(n3735), .ZN(n4476) );
  OAI22_X1 U4085 ( .A1(n3737), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[10][13] ), .B2(n3735), .ZN(n4477) );
  OAI22_X1 U4086 ( .A1(n3737), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[10][14] ), .B2(n3735), .ZN(n4478) );
  OAI22_X1 U4087 ( .A1(n3737), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[10][15] ), .B2(n3736), .ZN(n4479) );
  OAI22_X1 U4088 ( .A1(n3737), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[10][16] ), .B2(n3735), .ZN(n4480) );
  OAI22_X1 U4089 ( .A1(n3737), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[10][17] ), .B2(n3735), .ZN(n4481) );
  OAI22_X1 U4090 ( .A1(n3737), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[10][18] ), .B2(n3735), .ZN(n4482) );
  OAI22_X1 U4091 ( .A1(n3737), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[10][19] ), .B2(n3736), .ZN(n4483) );
  OAI22_X1 U4092 ( .A1(n3737), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[10][20] ), .B2(n3735), .ZN(n4484) );
  OAI22_X1 U4093 ( .A1(n3737), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[10][21] ), .B2(n3735), .ZN(n4485) );
  OAI22_X1 U4094 ( .A1(n3737), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[10][22] ), .B2(n3736), .ZN(n4486) );
  OAI22_X1 U4095 ( .A1(n3737), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[10][23] ), .B2(n3736), .ZN(n4487) );
  OAI22_X1 U4096 ( .A1(n3737), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[10][24] ), .B2(n3736), .ZN(n4488) );
  OAI22_X1 U4097 ( .A1(n3737), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[10][25] ), .B2(n3735), .ZN(n4489) );
  OAI22_X1 U4098 ( .A1(n3737), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[10][26] ), .B2(n3736), .ZN(n4490) );
  OAI22_X1 U4099 ( .A1(n3737), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[10][27] ), .B2(n3735), .ZN(n4491) );
  OAI22_X1 U4100 ( .A1(n3737), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[10][28] ), .B2(n3736), .ZN(n4492) );
  OAI22_X1 U4101 ( .A1(n3737), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[10][29] ), .B2(n3735), .ZN(n4493) );
  OAI22_X1 U4102 ( .A1(n3737), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[10][30] ), .B2(n3736), .ZN(n4494) );
  OAI22_X1 U4103 ( .A1(n3737), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[10][31] ), .B2(n3736), .ZN(n4495) );
  NOR2_X2 U4104 ( .A1(n3873), .A2(n3750), .ZN(n3738) );
  INV_X2 U4105 ( .A(n3739), .ZN(n3740) );
  OAI22_X1 U4106 ( .A1(n3740), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[11][0] ), .B2(n3739), .ZN(n4496) );
  OAI22_X1 U4107 ( .A1(n3740), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[11][1] ), .B2(n3738), .ZN(n4497) );
  OAI22_X1 U4108 ( .A1(n3740), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[11][2] ), .B2(n3738), .ZN(n4498) );
  OAI22_X1 U4109 ( .A1(n3740), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[11][3] ), .B2(n3738), .ZN(n4499) );
  OAI22_X1 U4110 ( .A1(n3740), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[11][4] ), .B2(n3738), .ZN(n4500) );
  OAI22_X1 U4111 ( .A1(n3740), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[11][5] ), .B2(n3738), .ZN(n4501) );
  OAI22_X1 U4112 ( .A1(n3740), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[11][6] ), .B2(n3738), .ZN(n4502) );
  OAI22_X1 U4113 ( .A1(n3740), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[11][7] ), .B2(n3738), .ZN(n4503) );
  OAI22_X1 U4114 ( .A1(n3740), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[11][8] ), .B2(n3738), .ZN(n4504) );
  OAI22_X1 U4115 ( .A1(n3740), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[11][9] ), .B2(n3738), .ZN(n4505) );
  OAI22_X1 U4116 ( .A1(n3740), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[11][10] ), .B2(n3738), .ZN(n4506) );
  OAI22_X1 U4117 ( .A1(n3740), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[11][11] ), .B2(n3738), .ZN(n4507) );
  OAI22_X1 U4118 ( .A1(n3740), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[11][12] ), .B2(n3738), .ZN(n4508) );
  OAI22_X1 U4119 ( .A1(n3740), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[11][13] ), .B2(n3738), .ZN(n4509) );
  OAI22_X1 U4120 ( .A1(n3740), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[11][14] ), .B2(n3738), .ZN(n4510) );
  OAI22_X1 U4121 ( .A1(n3740), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[11][15] ), .B2(n3739), .ZN(n4511) );
  OAI22_X1 U4122 ( .A1(n3740), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[11][16] ), .B2(n3738), .ZN(n4512) );
  OAI22_X1 U4123 ( .A1(n3740), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[11][17] ), .B2(n3738), .ZN(n4513) );
  OAI22_X1 U4124 ( .A1(n3740), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[11][18] ), .B2(n3738), .ZN(n4514) );
  OAI22_X1 U4125 ( .A1(n3740), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[11][19] ), .B2(n3739), .ZN(n4515) );
  OAI22_X1 U4126 ( .A1(n3740), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[11][20] ), .B2(n3738), .ZN(n4516) );
  OAI22_X1 U4127 ( .A1(n3740), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[11][21] ), .B2(n3738), .ZN(n4517) );
  OAI22_X1 U4128 ( .A1(n3740), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[11][22] ), .B2(n3739), .ZN(n4518) );
  OAI22_X1 U4129 ( .A1(n3740), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[11][23] ), .B2(n3739), .ZN(n4519) );
  OAI22_X1 U4130 ( .A1(n3740), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[11][24] ), .B2(n3739), .ZN(n4520) );
  OAI22_X1 U4131 ( .A1(n3740), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[11][25] ), .B2(n3738), .ZN(n4521) );
  OAI22_X1 U4132 ( .A1(n3740), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[11][26] ), .B2(n3739), .ZN(n4522) );
  OAI22_X1 U4133 ( .A1(n3740), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[11][27] ), .B2(n3738), .ZN(n4523) );
  OAI22_X1 U4134 ( .A1(n3740), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[11][28] ), .B2(n3739), .ZN(n4524) );
  OAI22_X1 U4135 ( .A1(n3740), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[11][29] ), .B2(n3738), .ZN(n4525) );
  OAI22_X1 U4136 ( .A1(n3740), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[11][30] ), .B2(n3739), .ZN(n4526) );
  OAI22_X1 U4137 ( .A1(n3740), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[11][31] ), .B2(n3739), .ZN(n4527) );
  NOR2_X2 U4138 ( .A1(n3878), .A2(n3750), .ZN(n3741) );
  INV_X2 U4139 ( .A(n3742), .ZN(n3743) );
  OAI22_X1 U4140 ( .A1(n3743), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[12][0] ), .B2(n3742), .ZN(n4528) );
  OAI22_X1 U4141 ( .A1(n3743), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[12][1] ), .B2(n3741), .ZN(n4529) );
  OAI22_X1 U4142 ( .A1(n3743), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[12][2] ), .B2(n3741), .ZN(n4530) );
  OAI22_X1 U4143 ( .A1(n3743), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[12][3] ), .B2(n3741), .ZN(n4531) );
  OAI22_X1 U4144 ( .A1(n3743), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[12][4] ), .B2(n3741), .ZN(n4532) );
  OAI22_X1 U4145 ( .A1(n3743), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[12][5] ), .B2(n3741), .ZN(n4533) );
  OAI22_X1 U4146 ( .A1(n3743), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[12][6] ), .B2(n3741), .ZN(n4534) );
  OAI22_X1 U4147 ( .A1(n3743), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[12][7] ), .B2(n3741), .ZN(n4535) );
  OAI22_X1 U4148 ( .A1(n3743), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[12][8] ), .B2(n3741), .ZN(n4536) );
  OAI22_X1 U4149 ( .A1(n3743), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[12][9] ), .B2(n3741), .ZN(n4537) );
  OAI22_X1 U4150 ( .A1(n3743), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[12][10] ), .B2(n3741), .ZN(n4538) );
  OAI22_X1 U4151 ( .A1(n3743), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[12][11] ), .B2(n3741), .ZN(n4539) );
  OAI22_X1 U4152 ( .A1(n3743), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[12][12] ), .B2(n3741), .ZN(n4540) );
  OAI22_X1 U4153 ( .A1(n3743), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[12][13] ), .B2(n3741), .ZN(n4541) );
  OAI22_X1 U4154 ( .A1(n3743), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[12][14] ), .B2(n3741), .ZN(n4542) );
  OAI22_X1 U4155 ( .A1(n3743), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[12][15] ), .B2(n3742), .ZN(n4543) );
  OAI22_X1 U4156 ( .A1(n3743), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[12][16] ), .B2(n3741), .ZN(n4544) );
  OAI22_X1 U4157 ( .A1(n3743), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[12][17] ), .B2(n3741), .ZN(n4545) );
  OAI22_X1 U4158 ( .A1(n3743), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[12][18] ), .B2(n3741), .ZN(n4546) );
  OAI22_X1 U4159 ( .A1(n3743), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[12][19] ), .B2(n3742), .ZN(n4547) );
  OAI22_X1 U4160 ( .A1(n3743), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[12][20] ), .B2(n3741), .ZN(n4548) );
  OAI22_X1 U4161 ( .A1(n3743), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[12][21] ), .B2(n3741), .ZN(n4549) );
  OAI22_X1 U4162 ( .A1(n3743), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[12][22] ), .B2(n3742), .ZN(n4550) );
  OAI22_X1 U4163 ( .A1(n3743), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[12][23] ), .B2(n3742), .ZN(n4551) );
  OAI22_X1 U4164 ( .A1(n3743), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[12][24] ), .B2(n3742), .ZN(n4552) );
  OAI22_X1 U4165 ( .A1(n3743), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[12][25] ), .B2(n3741), .ZN(n4553) );
  OAI22_X1 U4166 ( .A1(n3743), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[12][26] ), .B2(n3742), .ZN(n4554) );
  OAI22_X1 U4167 ( .A1(n3743), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[12][27] ), .B2(n3741), .ZN(n4555) );
  OAI22_X1 U4168 ( .A1(n3743), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[12][28] ), .B2(n3742), .ZN(n4556) );
  OAI22_X1 U4169 ( .A1(n3743), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[12][29] ), .B2(n3741), .ZN(n4557) );
  OAI22_X1 U4170 ( .A1(n3743), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[12][30] ), .B2(n3742), .ZN(n4558) );
  OAI22_X1 U4171 ( .A1(n3743), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[12][31] ), .B2(n3742), .ZN(n4559) );
  NOR2_X2 U4172 ( .A1(n3882), .A2(n3750), .ZN(n3744) );
  INV_X2 U4173 ( .A(n3745), .ZN(n3746) );
  OAI22_X1 U4174 ( .A1(n3746), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[13][0] ), .B2(n3745), .ZN(n4560) );
  OAI22_X1 U4175 ( .A1(n3746), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[13][1] ), .B2(n3744), .ZN(n4561) );
  OAI22_X1 U4176 ( .A1(n3746), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[13][2] ), .B2(n3744), .ZN(n4562) );
  OAI22_X1 U4177 ( .A1(n3746), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[13][3] ), .B2(n3744), .ZN(n4563) );
  OAI22_X1 U4178 ( .A1(n3746), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[13][4] ), .B2(n3744), .ZN(n4564) );
  OAI22_X1 U4179 ( .A1(n3746), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[13][5] ), .B2(n3744), .ZN(n4565) );
  OAI22_X1 U4180 ( .A1(n3746), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[13][6] ), .B2(n3744), .ZN(n4566) );
  OAI22_X1 U4181 ( .A1(n3746), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[13][7] ), .B2(n3744), .ZN(n4567) );
  OAI22_X1 U4182 ( .A1(n3746), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[13][8] ), .B2(n3744), .ZN(n4568) );
  OAI22_X1 U4183 ( .A1(n3746), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[13][9] ), .B2(n3744), .ZN(n4569) );
  OAI22_X1 U4184 ( .A1(n3746), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[13][10] ), .B2(n3744), .ZN(n4570) );
  OAI22_X1 U4185 ( .A1(n3746), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[13][11] ), .B2(n3744), .ZN(n4571) );
  OAI22_X1 U4186 ( .A1(n3746), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[13][12] ), .B2(n3744), .ZN(n4572) );
  OAI22_X1 U4187 ( .A1(n3746), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[13][13] ), .B2(n3744), .ZN(n4573) );
  OAI22_X1 U4188 ( .A1(n3746), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[13][14] ), .B2(n3744), .ZN(n4574) );
  OAI22_X1 U4189 ( .A1(n3746), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[13][15] ), .B2(n3745), .ZN(n4575) );
  OAI22_X1 U4190 ( .A1(n3746), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[13][16] ), .B2(n3744), .ZN(n4576) );
  OAI22_X1 U4191 ( .A1(n3746), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[13][17] ), .B2(n3744), .ZN(n4577) );
  OAI22_X1 U4192 ( .A1(n3746), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[13][18] ), .B2(n3744), .ZN(n4578) );
  OAI22_X1 U4193 ( .A1(n3746), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[13][19] ), .B2(n3745), .ZN(n4579) );
  OAI22_X1 U4194 ( .A1(n3746), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[13][20] ), .B2(n3744), .ZN(n4580) );
  OAI22_X1 U4195 ( .A1(n3746), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[13][21] ), .B2(n3744), .ZN(n4581) );
  OAI22_X1 U4196 ( .A1(n3746), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[13][22] ), .B2(n3745), .ZN(n4582) );
  OAI22_X1 U4197 ( .A1(n3746), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[13][23] ), .B2(n3745), .ZN(n4583) );
  OAI22_X1 U4198 ( .A1(n3746), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[13][24] ), .B2(n3745), .ZN(n4584) );
  OAI22_X1 U4199 ( .A1(n3746), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[13][25] ), .B2(n3744), .ZN(n4585) );
  OAI22_X1 U4200 ( .A1(n3746), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[13][26] ), .B2(n3745), .ZN(n4586) );
  OAI22_X1 U4201 ( .A1(n3746), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[13][27] ), .B2(n3744), .ZN(n4587) );
  OAI22_X1 U4202 ( .A1(n3746), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[13][28] ), .B2(n3745), .ZN(n4588) );
  OAI22_X1 U4203 ( .A1(n3746), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[13][29] ), .B2(n3744), .ZN(n4589) );
  OAI22_X1 U4204 ( .A1(n3746), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[13][30] ), .B2(n3745), .ZN(n4590) );
  OAI22_X1 U4205 ( .A1(n3746), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[13][31] ), .B2(n3745), .ZN(n4591) );
  NOR2_X2 U4206 ( .A1(n3886), .A2(n3750), .ZN(n3747) );
  INV_X2 U4207 ( .A(n3748), .ZN(n3749) );
  OAI22_X1 U4208 ( .A1(n3749), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[14][0] ), .B2(n3748), .ZN(n4592) );
  OAI22_X1 U4209 ( .A1(n3749), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[14][1] ), .B2(n3747), .ZN(n4593) );
  OAI22_X1 U4210 ( .A1(n3749), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[14][2] ), .B2(n3747), .ZN(n4594) );
  OAI22_X1 U4211 ( .A1(n3749), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[14][3] ), .B2(n3747), .ZN(n4595) );
  OAI22_X1 U4212 ( .A1(n3749), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[14][4] ), .B2(n3747), .ZN(n4596) );
  OAI22_X1 U4213 ( .A1(n3749), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[14][5] ), .B2(n3747), .ZN(n4597) );
  OAI22_X1 U4214 ( .A1(n3749), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[14][6] ), .B2(n3747), .ZN(n4598) );
  OAI22_X1 U4215 ( .A1(n3749), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[14][7] ), .B2(n3747), .ZN(n4599) );
  OAI22_X1 U4216 ( .A1(n3749), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[14][8] ), .B2(n3747), .ZN(n4600) );
  OAI22_X1 U4217 ( .A1(n3749), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[14][9] ), .B2(n3747), .ZN(n4601) );
  OAI22_X1 U4218 ( .A1(n3749), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[14][10] ), .B2(n3747), .ZN(n4602) );
  OAI22_X1 U4219 ( .A1(n3749), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[14][11] ), .B2(n3747), .ZN(n4603) );
  OAI22_X1 U4220 ( .A1(n3749), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[14][12] ), .B2(n3747), .ZN(n4604) );
  OAI22_X1 U4221 ( .A1(n3749), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[14][13] ), .B2(n3747), .ZN(n4605) );
  OAI22_X1 U4222 ( .A1(n3749), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[14][14] ), .B2(n3747), .ZN(n4606) );
  OAI22_X1 U4223 ( .A1(n3749), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[14][15] ), .B2(n3748), .ZN(n4607) );
  OAI22_X1 U4224 ( .A1(n3749), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[14][16] ), .B2(n3747), .ZN(n4608) );
  OAI22_X1 U4225 ( .A1(n3749), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[14][17] ), .B2(n3747), .ZN(n4609) );
  OAI22_X1 U4226 ( .A1(n3749), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[14][18] ), .B2(n3747), .ZN(n4610) );
  OAI22_X1 U4227 ( .A1(n3749), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[14][19] ), .B2(n3748), .ZN(n4611) );
  OAI22_X1 U4228 ( .A1(n3749), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[14][20] ), .B2(n3747), .ZN(n4612) );
  OAI22_X1 U4229 ( .A1(n3749), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[14][21] ), .B2(n3747), .ZN(n4613) );
  OAI22_X1 U4230 ( .A1(n3749), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[14][22] ), .B2(n3748), .ZN(n4614) );
  OAI22_X1 U4231 ( .A1(n3749), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[14][23] ), .B2(n3748), .ZN(n4615) );
  OAI22_X1 U4232 ( .A1(n3749), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[14][24] ), .B2(n3748), .ZN(n4616) );
  OAI22_X1 U4233 ( .A1(n3749), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[14][25] ), .B2(n3747), .ZN(n4617) );
  OAI22_X1 U4234 ( .A1(n3749), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[14][26] ), .B2(n3748), .ZN(n4618) );
  OAI22_X1 U4235 ( .A1(n3749), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[14][27] ), .B2(n3747), .ZN(n4619) );
  OAI22_X1 U4236 ( .A1(n3749), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[14][28] ), .B2(n3748), .ZN(n4620) );
  OAI22_X1 U4237 ( .A1(n3749), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[14][29] ), .B2(n3747), .ZN(n4621) );
  OAI22_X1 U4238 ( .A1(n3749), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[14][30] ), .B2(n3748), .ZN(n4622) );
  OAI22_X1 U4239 ( .A1(n3749), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[14][31] ), .B2(n3748), .ZN(n4623) );
  NOR2_X2 U4240 ( .A1(n3891), .A2(n3750), .ZN(n3751) );
  INV_X2 U4241 ( .A(n3752), .ZN(n3753) );
  OAI22_X1 U4242 ( .A1(n3753), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[15][0] ), .B2(n3752), .ZN(n4624) );
  OAI22_X1 U4243 ( .A1(n3753), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[15][1] ), .B2(n3751), .ZN(n4625) );
  OAI22_X1 U4244 ( .A1(n3753), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[15][2] ), .B2(n3751), .ZN(n4626) );
  OAI22_X1 U4245 ( .A1(n3753), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[15][3] ), .B2(n3751), .ZN(n4627) );
  OAI22_X1 U4246 ( .A1(n3753), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[15][4] ), .B2(n3751), .ZN(n4628) );
  OAI22_X1 U4247 ( .A1(n3753), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[15][5] ), .B2(n3751), .ZN(n4629) );
  OAI22_X1 U4248 ( .A1(n3753), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[15][6] ), .B2(n3751), .ZN(n4630) );
  OAI22_X1 U4249 ( .A1(n3753), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[15][7] ), .B2(n3751), .ZN(n4631) );
  OAI22_X1 U4250 ( .A1(n3753), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[15][8] ), .B2(n3751), .ZN(n4632) );
  OAI22_X1 U4251 ( .A1(n3753), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[15][9] ), .B2(n3751), .ZN(n4633) );
  OAI22_X1 U4252 ( .A1(n3753), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[15][10] ), .B2(n3751), .ZN(n4634) );
  OAI22_X1 U4253 ( .A1(n3753), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[15][11] ), .B2(n3751), .ZN(n4635) );
  OAI22_X1 U4254 ( .A1(n3753), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[15][12] ), .B2(n3751), .ZN(n4636) );
  OAI22_X1 U4255 ( .A1(n3753), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[15][13] ), .B2(n3751), .ZN(n4637) );
  OAI22_X1 U4256 ( .A1(n3753), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[15][14] ), .B2(n3751), .ZN(n4638) );
  OAI22_X1 U4257 ( .A1(n3753), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[15][15] ), .B2(n3752), .ZN(n4639) );
  OAI22_X1 U4258 ( .A1(n3753), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[15][16] ), .B2(n3751), .ZN(n4640) );
  OAI22_X1 U4259 ( .A1(n3753), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[15][17] ), .B2(n3751), .ZN(n4641) );
  OAI22_X1 U4260 ( .A1(n3753), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[15][18] ), .B2(n3751), .ZN(n4642) );
  OAI22_X1 U4261 ( .A1(n3753), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[15][19] ), .B2(n3752), .ZN(n4643) );
  OAI22_X1 U4262 ( .A1(n3753), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[15][20] ), .B2(n3751), .ZN(n4644) );
  OAI22_X1 U4263 ( .A1(n3753), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[15][21] ), .B2(n3751), .ZN(n4645) );
  OAI22_X1 U4264 ( .A1(n3753), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[15][22] ), .B2(n3752), .ZN(n4646) );
  OAI22_X1 U4265 ( .A1(n3753), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[15][23] ), .B2(n3752), .ZN(n4647) );
  OAI22_X1 U4266 ( .A1(n3753), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[15][24] ), .B2(n3752), .ZN(n4648) );
  OAI22_X1 U4267 ( .A1(n3753), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[15][25] ), .B2(n3751), .ZN(n4649) );
  OAI22_X1 U4268 ( .A1(n3753), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[15][26] ), .B2(n3752), .ZN(n4650) );
  OAI22_X1 U4269 ( .A1(n3753), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[15][27] ), .B2(n3751), .ZN(n4651) );
  OAI22_X1 U4270 ( .A1(n3753), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[15][28] ), .B2(n3752), .ZN(n4652) );
  OAI22_X1 U4271 ( .A1(n3753), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[15][29] ), .B2(n3751), .ZN(n4653) );
  OAI22_X1 U4272 ( .A1(n3753), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[15][30] ), .B2(n3752), .ZN(n4654) );
  OAI22_X1 U4273 ( .A1(n3753), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[15][31] ), .B2(n3752), .ZN(n4655) );
  NOR2_X2 U4274 ( .A1(n3897), .A2(n3775), .ZN(n3754) );
  INV_X2 U4275 ( .A(n3755), .ZN(n3756) );
  OAI22_X1 U4276 ( .A1(n3756), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[16][0] ), .B2(n3755), .ZN(n4656) );
  OAI22_X1 U4277 ( .A1(n3756), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[16][1] ), .B2(n3754), .ZN(n4657) );
  OAI22_X1 U4278 ( .A1(n3756), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[16][2] ), .B2(n3754), .ZN(n4658) );
  OAI22_X1 U4279 ( .A1(n3756), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[16][3] ), .B2(n3754), .ZN(n4659) );
  OAI22_X1 U4280 ( .A1(n3756), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[16][4] ), .B2(n3754), .ZN(n4660) );
  OAI22_X1 U4281 ( .A1(n3756), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[16][5] ), .B2(n3754), .ZN(n4661) );
  OAI22_X1 U4282 ( .A1(n3756), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[16][6] ), .B2(n3754), .ZN(n4662) );
  OAI22_X1 U4283 ( .A1(n3756), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[16][7] ), .B2(n3754), .ZN(n4663) );
  OAI22_X1 U4284 ( .A1(n3756), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[16][8] ), .B2(n3754), .ZN(n4664) );
  OAI22_X1 U4285 ( .A1(n3756), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[16][9] ), .B2(n3754), .ZN(n4665) );
  OAI22_X1 U4286 ( .A1(n3756), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[16][10] ), .B2(n3754), .ZN(n4666) );
  OAI22_X1 U4287 ( .A1(n3756), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[16][11] ), .B2(n3754), .ZN(n4667) );
  OAI22_X1 U4288 ( .A1(n3756), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[16][12] ), .B2(n3754), .ZN(n4668) );
  OAI22_X1 U4289 ( .A1(n3756), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[16][13] ), .B2(n3754), .ZN(n4669) );
  OAI22_X1 U4290 ( .A1(n3756), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[16][14] ), .B2(n3754), .ZN(n4670) );
  OAI22_X1 U4291 ( .A1(n3756), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[16][15] ), .B2(n3755), .ZN(n4671) );
  OAI22_X1 U4292 ( .A1(n3756), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[16][16] ), .B2(n3754), .ZN(n4672) );
  OAI22_X1 U4293 ( .A1(n3756), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[16][17] ), .B2(n3754), .ZN(n4673) );
  OAI22_X1 U4294 ( .A1(n3756), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[16][18] ), .B2(n3754), .ZN(n4674) );
  OAI22_X1 U4295 ( .A1(n3756), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[16][19] ), .B2(n3755), .ZN(n4675) );
  OAI22_X1 U4296 ( .A1(n3756), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[16][20] ), .B2(n3754), .ZN(n4676) );
  OAI22_X1 U4297 ( .A1(n3756), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[16][21] ), .B2(n3754), .ZN(n4677) );
  OAI22_X1 U4298 ( .A1(n3756), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[16][22] ), .B2(n3755), .ZN(n4678) );
  OAI22_X1 U4299 ( .A1(n3756), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[16][23] ), .B2(n3755), .ZN(n4679) );
  OAI22_X1 U4300 ( .A1(n3756), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[16][24] ), .B2(n3755), .ZN(n4680) );
  OAI22_X1 U4301 ( .A1(n3756), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[16][25] ), .B2(n3754), .ZN(n4681) );
  OAI22_X1 U4302 ( .A1(n3756), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[16][26] ), .B2(n3755), .ZN(n4682) );
  OAI22_X1 U4303 ( .A1(n3756), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[16][27] ), .B2(n3754), .ZN(n4683) );
  OAI22_X1 U4304 ( .A1(n3756), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[16][28] ), .B2(n3755), .ZN(n4684) );
  OAI22_X1 U4305 ( .A1(n3756), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[16][29] ), .B2(n3754), .ZN(n4685) );
  OAI22_X1 U4306 ( .A1(n3756), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[16][30] ), .B2(n3755), .ZN(n4686) );
  OAI22_X1 U4307 ( .A1(n3756), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[16][31] ), .B2(n3755), .ZN(n4687) );
  NOR2_X2 U4308 ( .A1(n3933), .A2(n3775), .ZN(n3757) );
  INV_X2 U4309 ( .A(n3758), .ZN(n3759) );
  OAI22_X1 U4310 ( .A1(n3759), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[17][0] ), .B2(n3758), .ZN(n4688) );
  OAI22_X1 U4311 ( .A1(n3759), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[17][1] ), .B2(n3757), .ZN(n4689) );
  OAI22_X1 U4312 ( .A1(n3759), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[17][2] ), .B2(n3757), .ZN(n4690) );
  OAI22_X1 U4313 ( .A1(n3759), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[17][3] ), .B2(n3757), .ZN(n4691) );
  OAI22_X1 U4314 ( .A1(n3759), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[17][4] ), .B2(n3757), .ZN(n4692) );
  OAI22_X1 U4315 ( .A1(n3759), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[17][5] ), .B2(n3757), .ZN(n4693) );
  OAI22_X1 U4316 ( .A1(n3759), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[17][6] ), .B2(n3757), .ZN(n4694) );
  OAI22_X1 U4317 ( .A1(n3759), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[17][7] ), .B2(n3757), .ZN(n4695) );
  OAI22_X1 U4318 ( .A1(n3759), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[17][8] ), .B2(n3757), .ZN(n4696) );
  OAI22_X1 U4319 ( .A1(n3759), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[17][9] ), .B2(n3757), .ZN(n4697) );
  OAI22_X1 U4320 ( .A1(n3759), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[17][10] ), .B2(n3757), .ZN(n4698) );
  OAI22_X1 U4321 ( .A1(n3759), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[17][11] ), .B2(n3757), .ZN(n4699) );
  OAI22_X1 U4322 ( .A1(n3759), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[17][12] ), .B2(n3757), .ZN(n4700) );
  OAI22_X1 U4323 ( .A1(n3759), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[17][13] ), .B2(n3757), .ZN(n4701) );
  OAI22_X1 U4324 ( .A1(n3759), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[17][14] ), .B2(n3757), .ZN(n4702) );
  OAI22_X1 U4325 ( .A1(n3759), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[17][15] ), .B2(n3758), .ZN(n4703) );
  OAI22_X1 U4326 ( .A1(n3759), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[17][16] ), .B2(n3757), .ZN(n4704) );
  OAI22_X1 U4327 ( .A1(n3759), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[17][17] ), .B2(n3757), .ZN(n4705) );
  OAI22_X1 U4328 ( .A1(n3759), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[17][18] ), .B2(n3757), .ZN(n4706) );
  OAI22_X1 U4329 ( .A1(n3759), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[17][19] ), .B2(n3758), .ZN(n4707) );
  OAI22_X1 U4330 ( .A1(n3759), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[17][20] ), .B2(n3757), .ZN(n4708) );
  OAI22_X1 U4331 ( .A1(n3759), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[17][21] ), .B2(n3757), .ZN(n4709) );
  OAI22_X1 U4332 ( .A1(n3759), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[17][22] ), .B2(n3758), .ZN(n4710) );
  OAI22_X1 U4333 ( .A1(n3759), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[17][23] ), .B2(n3758), .ZN(n4711) );
  OAI22_X1 U4334 ( .A1(n3759), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[17][24] ), .B2(n3758), .ZN(n4712) );
  OAI22_X1 U4335 ( .A1(n3759), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[17][25] ), .B2(n3757), .ZN(n4713) );
  OAI22_X1 U4336 ( .A1(n3759), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[17][26] ), .B2(n3758), .ZN(n4714) );
  OAI22_X1 U4337 ( .A1(n3759), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[17][27] ), .B2(n3757), .ZN(n4715) );
  OAI22_X1 U4338 ( .A1(n3759), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[17][28] ), .B2(n3758), .ZN(n4716) );
  OAI22_X1 U4339 ( .A1(n3759), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[17][29] ), .B2(n3757), .ZN(n4717) );
  OAI22_X1 U4340 ( .A1(n3759), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[17][30] ), .B2(n3758), .ZN(n4718) );
  OAI22_X1 U4341 ( .A1(n3759), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[17][31] ), .B2(n3758), .ZN(n4719) );
  NOR2_X2 U4342 ( .A1(n3970), .A2(n3775), .ZN(n3760) );
  INV_X2 U4343 ( .A(n3761), .ZN(n3762) );
  OAI22_X1 U4344 ( .A1(n3762), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[18][0] ), .B2(n3761), .ZN(n4720) );
  OAI22_X1 U4345 ( .A1(n3762), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[18][1] ), .B2(n3760), .ZN(n4721) );
  OAI22_X1 U4346 ( .A1(n3762), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[18][2] ), .B2(n3760), .ZN(n4722) );
  OAI22_X1 U4347 ( .A1(n3762), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[18][3] ), .B2(n3760), .ZN(n4723) );
  OAI22_X1 U4348 ( .A1(n3762), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[18][4] ), .B2(n3760), .ZN(n4724) );
  OAI22_X1 U4349 ( .A1(n3762), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[18][5] ), .B2(n3760), .ZN(n4725) );
  OAI22_X1 U4350 ( .A1(n3762), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[18][6] ), .B2(n3760), .ZN(n4726) );
  OAI22_X1 U4351 ( .A1(n3762), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[18][7] ), .B2(n3760), .ZN(n4727) );
  OAI22_X1 U4352 ( .A1(n3762), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[18][8] ), .B2(n3760), .ZN(n4728) );
  OAI22_X1 U4353 ( .A1(n3762), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[18][9] ), .B2(n3760), .ZN(n4729) );
  OAI22_X1 U4354 ( .A1(n3762), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[18][10] ), .B2(n3760), .ZN(n4730) );
  OAI22_X1 U4355 ( .A1(n3762), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[18][11] ), .B2(n3760), .ZN(n4731) );
  OAI22_X1 U4356 ( .A1(n3762), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[18][12] ), .B2(n3760), .ZN(n4732) );
  OAI22_X1 U4357 ( .A1(n3762), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[18][13] ), .B2(n3760), .ZN(n4733) );
  OAI22_X1 U4358 ( .A1(n3762), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[18][14] ), .B2(n3760), .ZN(n4734) );
  OAI22_X1 U4359 ( .A1(n3762), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[18][15] ), .B2(n3761), .ZN(n4735) );
  OAI22_X1 U4360 ( .A1(n3762), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[18][16] ), .B2(n3760), .ZN(n4736) );
  OAI22_X1 U4361 ( .A1(n3762), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[18][17] ), .B2(n3760), .ZN(n4737) );
  OAI22_X1 U4362 ( .A1(n3762), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[18][18] ), .B2(n3760), .ZN(n4738) );
  OAI22_X1 U4363 ( .A1(n3762), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[18][19] ), .B2(n3761), .ZN(n4739) );
  OAI22_X1 U4364 ( .A1(n3762), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[18][20] ), .B2(n3760), .ZN(n4740) );
  OAI22_X1 U4365 ( .A1(n3762), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[18][21] ), .B2(n3760), .ZN(n4741) );
  OAI22_X1 U4366 ( .A1(n3762), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[18][22] ), .B2(n3761), .ZN(n4742) );
  OAI22_X1 U4367 ( .A1(n3762), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[18][23] ), .B2(n3761), .ZN(n4743) );
  OAI22_X1 U4368 ( .A1(n3762), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[18][24] ), .B2(n3761), .ZN(n4744) );
  OAI22_X1 U4369 ( .A1(n3762), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[18][25] ), .B2(n3760), .ZN(n4745) );
  OAI22_X1 U4370 ( .A1(n3762), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[18][26] ), .B2(n3761), .ZN(n4746) );
  OAI22_X1 U4371 ( .A1(n3762), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[18][27] ), .B2(n3760), .ZN(n4747) );
  OAI22_X1 U4372 ( .A1(n3762), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[18][28] ), .B2(n3761), .ZN(n4748) );
  OAI22_X1 U4373 ( .A1(n3762), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[18][29] ), .B2(n3760), .ZN(n4749) );
  OAI22_X1 U4374 ( .A1(n3762), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[18][30] ), .B2(n3761), .ZN(n4750) );
  OAI22_X1 U4375 ( .A1(n3762), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[18][31] ), .B2(n3761), .ZN(n4751) );
  NOR2_X2 U4376 ( .A1(n3873), .A2(n3775), .ZN(n3763) );
  INV_X2 U4377 ( .A(n3764), .ZN(n3765) );
  OAI22_X1 U4378 ( .A1(n3765), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[19][0] ), .B2(n3764), .ZN(n4752) );
  OAI22_X1 U4379 ( .A1(n3765), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[19][1] ), .B2(n3763), .ZN(n4753) );
  OAI22_X1 U4380 ( .A1(n3765), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[19][2] ), .B2(n3763), .ZN(n4754) );
  OAI22_X1 U4381 ( .A1(n3765), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[19][3] ), .B2(n3763), .ZN(n4755) );
  OAI22_X1 U4382 ( .A1(n3765), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[19][4] ), .B2(n3763), .ZN(n4756) );
  OAI22_X1 U4383 ( .A1(n3765), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[19][5] ), .B2(n3763), .ZN(n4757) );
  OAI22_X1 U4384 ( .A1(n3765), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[19][6] ), .B2(n3763), .ZN(n4758) );
  OAI22_X1 U4385 ( .A1(n3765), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[19][7] ), .B2(n3763), .ZN(n4759) );
  OAI22_X1 U4386 ( .A1(n3765), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[19][8] ), .B2(n3763), .ZN(n4760) );
  OAI22_X1 U4387 ( .A1(n3765), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[19][9] ), .B2(n3763), .ZN(n4761) );
  OAI22_X1 U4388 ( .A1(n3765), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[19][10] ), .B2(n3763), .ZN(n4762) );
  OAI22_X1 U4389 ( .A1(n3765), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[19][11] ), .B2(n3763), .ZN(n4763) );
  OAI22_X1 U4390 ( .A1(n3765), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[19][12] ), .B2(n3763), .ZN(n4764) );
  OAI22_X1 U4391 ( .A1(n3765), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[19][13] ), .B2(n3763), .ZN(n4765) );
  OAI22_X1 U4392 ( .A1(n3765), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[19][14] ), .B2(n3763), .ZN(n4766) );
  OAI22_X1 U4393 ( .A1(n3765), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[19][15] ), .B2(n3764), .ZN(n4767) );
  OAI22_X1 U4394 ( .A1(n3765), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[19][16] ), .B2(n3763), .ZN(n4768) );
  OAI22_X1 U4395 ( .A1(n3765), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[19][17] ), .B2(n3763), .ZN(n4769) );
  OAI22_X1 U4396 ( .A1(n3765), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[19][18] ), .B2(n3763), .ZN(n4770) );
  OAI22_X1 U4397 ( .A1(n3765), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[19][19] ), .B2(n3764), .ZN(n4771) );
  OAI22_X1 U4398 ( .A1(n3765), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[19][20] ), .B2(n3763), .ZN(n4772) );
  OAI22_X1 U4399 ( .A1(n3765), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[19][21] ), .B2(n3763), .ZN(n4773) );
  OAI22_X1 U4400 ( .A1(n3765), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[19][22] ), .B2(n3764), .ZN(n4774) );
  OAI22_X1 U4401 ( .A1(n3765), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[19][23] ), .B2(n3764), .ZN(n4775) );
  OAI22_X1 U4402 ( .A1(n3765), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[19][24] ), .B2(n3764), .ZN(n4776) );
  OAI22_X1 U4403 ( .A1(n3765), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[19][25] ), .B2(n3763), .ZN(n4777) );
  OAI22_X1 U4404 ( .A1(n3765), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[19][26] ), .B2(n3764), .ZN(n4778) );
  OAI22_X1 U4405 ( .A1(n3765), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[19][27] ), .B2(n3763), .ZN(n4779) );
  OAI22_X1 U4406 ( .A1(n3765), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[19][28] ), .B2(n3764), .ZN(n4780) );
  OAI22_X1 U4407 ( .A1(n3765), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[19][29] ), .B2(n3763), .ZN(n4781) );
  OAI22_X1 U4408 ( .A1(n3765), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[19][30] ), .B2(n3764), .ZN(n4782) );
  OAI22_X1 U4409 ( .A1(n3765), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[19][31] ), .B2(n3764), .ZN(n4783) );
  NOR2_X2 U4410 ( .A1(n3878), .A2(n3775), .ZN(n3766) );
  INV_X2 U4411 ( .A(n3767), .ZN(n3768) );
  OAI22_X1 U4412 ( .A1(n3768), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[20][0] ), .B2(n3767), .ZN(n4784) );
  OAI22_X1 U4413 ( .A1(n3768), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[20][1] ), .B2(n3766), .ZN(n4785) );
  OAI22_X1 U4414 ( .A1(n3768), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[20][2] ), .B2(n3766), .ZN(n4786) );
  OAI22_X1 U4415 ( .A1(n3768), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[20][3] ), .B2(n3766), .ZN(n4787) );
  OAI22_X1 U4416 ( .A1(n3768), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[20][4] ), .B2(n3766), .ZN(n4788) );
  OAI22_X1 U4417 ( .A1(n3768), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[20][5] ), .B2(n3766), .ZN(n4789) );
  OAI22_X1 U4418 ( .A1(n3768), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[20][6] ), .B2(n3766), .ZN(n4790) );
  OAI22_X1 U4419 ( .A1(n3768), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[20][7] ), .B2(n3766), .ZN(n4791) );
  OAI22_X1 U4420 ( .A1(n3768), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[20][8] ), .B2(n3766), .ZN(n4792) );
  OAI22_X1 U4421 ( .A1(n3768), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[20][9] ), .B2(n3766), .ZN(n4793) );
  OAI22_X1 U4422 ( .A1(n3768), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[20][10] ), .B2(n3766), .ZN(n4794) );
  OAI22_X1 U4423 ( .A1(n3768), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[20][11] ), .B2(n3766), .ZN(n4795) );
  OAI22_X1 U4424 ( .A1(n3768), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[20][12] ), .B2(n3766), .ZN(n4796) );
  OAI22_X1 U4425 ( .A1(n3768), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[20][13] ), .B2(n3766), .ZN(n4797) );
  OAI22_X1 U4426 ( .A1(n3768), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[20][14] ), .B2(n3766), .ZN(n4798) );
  OAI22_X1 U4427 ( .A1(n3768), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[20][15] ), .B2(n3767), .ZN(n4799) );
  OAI22_X1 U4428 ( .A1(n3768), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[20][16] ), .B2(n3766), .ZN(n4800) );
  OAI22_X1 U4429 ( .A1(n3768), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[20][17] ), .B2(n3766), .ZN(n4801) );
  OAI22_X1 U4430 ( .A1(n3768), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[20][18] ), .B2(n3766), .ZN(n4802) );
  OAI22_X1 U4431 ( .A1(n3768), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[20][19] ), .B2(n3767), .ZN(n4803) );
  OAI22_X1 U4432 ( .A1(n3768), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[20][20] ), .B2(n3766), .ZN(n4804) );
  OAI22_X1 U4433 ( .A1(n3768), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[20][21] ), .B2(n3766), .ZN(n4805) );
  OAI22_X1 U4434 ( .A1(n3768), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[20][22] ), .B2(n3767), .ZN(n4806) );
  OAI22_X1 U4435 ( .A1(n3768), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[20][23] ), .B2(n3767), .ZN(n4807) );
  OAI22_X1 U4436 ( .A1(n3768), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[20][24] ), .B2(n3767), .ZN(n4808) );
  OAI22_X1 U4437 ( .A1(n3768), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[20][25] ), .B2(n3766), .ZN(n4809) );
  OAI22_X1 U4438 ( .A1(n3768), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[20][26] ), .B2(n3767), .ZN(n4810) );
  OAI22_X1 U4439 ( .A1(n3768), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[20][27] ), .B2(n3766), .ZN(n4811) );
  OAI22_X1 U4440 ( .A1(n3768), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[20][28] ), .B2(n3767), .ZN(n4812) );
  OAI22_X1 U4441 ( .A1(n3768), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[20][29] ), .B2(n3766), .ZN(n4813) );
  OAI22_X1 U4442 ( .A1(n3768), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[20][30] ), .B2(n3767), .ZN(n4814) );
  OAI22_X1 U4443 ( .A1(n3768), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[20][31] ), .B2(n3767), .ZN(n4815) );
  NOR2_X2 U4444 ( .A1(n3882), .A2(n3775), .ZN(n3769) );
  INV_X2 U4445 ( .A(n3770), .ZN(n3771) );
  OAI22_X1 U4446 ( .A1(n3771), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[21][0] ), .B2(n3770), .ZN(n4816) );
  OAI22_X1 U4447 ( .A1(n3771), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[21][1] ), .B2(n3769), .ZN(n4817) );
  OAI22_X1 U4448 ( .A1(n3771), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[21][2] ), .B2(n3769), .ZN(n4818) );
  OAI22_X1 U4449 ( .A1(n3771), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[21][3] ), .B2(n3769), .ZN(n4819) );
  OAI22_X1 U4450 ( .A1(n3771), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[21][4] ), .B2(n3769), .ZN(n4820) );
  OAI22_X1 U4451 ( .A1(n3771), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[21][5] ), .B2(n3769), .ZN(n4821) );
  OAI22_X1 U4452 ( .A1(n3771), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[21][6] ), .B2(n3769), .ZN(n4822) );
  OAI22_X1 U4453 ( .A1(n3771), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[21][7] ), .B2(n3769), .ZN(n4823) );
  OAI22_X1 U4454 ( .A1(n3771), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[21][8] ), .B2(n3769), .ZN(n4824) );
  OAI22_X1 U4455 ( .A1(n3771), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[21][9] ), .B2(n3769), .ZN(n4825) );
  OAI22_X1 U4456 ( .A1(n3771), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[21][10] ), .B2(n3769), .ZN(n4826) );
  OAI22_X1 U4457 ( .A1(n3771), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[21][11] ), .B2(n3769), .ZN(n4827) );
  OAI22_X1 U4458 ( .A1(n3771), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[21][12] ), .B2(n3769), .ZN(n4828) );
  OAI22_X1 U4459 ( .A1(n3771), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[21][13] ), .B2(n3769), .ZN(n4829) );
  OAI22_X1 U4460 ( .A1(n3771), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[21][14] ), .B2(n3769), .ZN(n4830) );
  OAI22_X1 U4461 ( .A1(n3771), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[21][15] ), .B2(n3770), .ZN(n4831) );
  OAI22_X1 U4462 ( .A1(n3771), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[21][16] ), .B2(n3769), .ZN(n4832) );
  OAI22_X1 U4463 ( .A1(n3771), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[21][17] ), .B2(n3769), .ZN(n4833) );
  OAI22_X1 U4464 ( .A1(n3771), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[21][18] ), .B2(n3769), .ZN(n4834) );
  OAI22_X1 U4465 ( .A1(n3771), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[21][19] ), .B2(n3770), .ZN(n4835) );
  OAI22_X1 U4466 ( .A1(n3771), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[21][20] ), .B2(n3769), .ZN(n4836) );
  OAI22_X1 U4467 ( .A1(n3771), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[21][21] ), .B2(n3769), .ZN(n4837) );
  OAI22_X1 U4468 ( .A1(n3771), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[21][22] ), .B2(n3770), .ZN(n4838) );
  OAI22_X1 U4469 ( .A1(n3771), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[21][23] ), .B2(n3770), .ZN(n4839) );
  OAI22_X1 U4470 ( .A1(n3771), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[21][24] ), .B2(n3770), .ZN(n4840) );
  OAI22_X1 U4471 ( .A1(n3771), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[21][25] ), .B2(n3769), .ZN(n4841) );
  OAI22_X1 U4472 ( .A1(n3771), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[21][26] ), .B2(n3770), .ZN(n4842) );
  OAI22_X1 U4473 ( .A1(n3771), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[21][27] ), .B2(n3769), .ZN(n4843) );
  OAI22_X1 U4474 ( .A1(n3771), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[21][28] ), .B2(n3770), .ZN(n4844) );
  OAI22_X1 U4475 ( .A1(n3771), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[21][29] ), .B2(n3769), .ZN(n4845) );
  OAI22_X1 U4476 ( .A1(n3771), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[21][30] ), .B2(n3770), .ZN(n4846) );
  OAI22_X1 U4477 ( .A1(n3771), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[21][31] ), .B2(n3770), .ZN(n4847) );
  NOR2_X2 U4478 ( .A1(n3886), .A2(n3775), .ZN(n3772) );
  INV_X2 U4479 ( .A(n3773), .ZN(n3774) );
  OAI22_X1 U4480 ( .A1(n3774), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[22][0] ), .B2(n3773), .ZN(n4848) );
  OAI22_X1 U4481 ( .A1(n3774), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[22][1] ), .B2(n3772), .ZN(n4849) );
  OAI22_X1 U4482 ( .A1(n3774), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[22][2] ), .B2(n3772), .ZN(n4850) );
  OAI22_X1 U4483 ( .A1(n3774), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[22][3] ), .B2(n3772), .ZN(n4851) );
  OAI22_X1 U4484 ( .A1(n3774), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[22][4] ), .B2(n3772), .ZN(n4852) );
  OAI22_X1 U4485 ( .A1(n3774), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[22][5] ), .B2(n3772), .ZN(n4853) );
  OAI22_X1 U4486 ( .A1(n3774), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[22][6] ), .B2(n3772), .ZN(n4854) );
  OAI22_X1 U4487 ( .A1(n3774), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[22][7] ), .B2(n3772), .ZN(n4855) );
  OAI22_X1 U4488 ( .A1(n3774), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[22][8] ), .B2(n3772), .ZN(n4856) );
  OAI22_X1 U4489 ( .A1(n3774), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[22][9] ), .B2(n3772), .ZN(n4857) );
  OAI22_X1 U4490 ( .A1(n3774), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[22][10] ), .B2(n3772), .ZN(n4858) );
  OAI22_X1 U4491 ( .A1(n3774), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[22][11] ), .B2(n3772), .ZN(n4859) );
  OAI22_X1 U4492 ( .A1(n3774), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[22][12] ), .B2(n3772), .ZN(n4860) );
  OAI22_X1 U4493 ( .A1(n3774), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[22][13] ), .B2(n3772), .ZN(n4861) );
  OAI22_X1 U4494 ( .A1(n3774), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[22][14] ), .B2(n3772), .ZN(n4862) );
  OAI22_X1 U4495 ( .A1(n3774), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[22][15] ), .B2(n3773), .ZN(n4863) );
  OAI22_X1 U4496 ( .A1(n3774), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[22][16] ), .B2(n3772), .ZN(n4864) );
  OAI22_X1 U4497 ( .A1(n3774), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[22][17] ), .B2(n3772), .ZN(n4865) );
  OAI22_X1 U4498 ( .A1(n3774), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[22][18] ), .B2(n3772), .ZN(n4866) );
  OAI22_X1 U4499 ( .A1(n3774), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[22][19] ), .B2(n3773), .ZN(n4867) );
  OAI22_X1 U4500 ( .A1(n3774), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[22][20] ), .B2(n3772), .ZN(n4868) );
  OAI22_X1 U4501 ( .A1(n3774), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[22][21] ), .B2(n3772), .ZN(n4869) );
  OAI22_X1 U4502 ( .A1(n3774), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[22][22] ), .B2(n3773), .ZN(n4870) );
  OAI22_X1 U4503 ( .A1(n3774), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[22][23] ), .B2(n3773), .ZN(n4871) );
  OAI22_X1 U4504 ( .A1(n3774), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[22][24] ), .B2(n3773), .ZN(n4872) );
  OAI22_X1 U4505 ( .A1(n3774), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[22][25] ), .B2(n3772), .ZN(n4873) );
  OAI22_X1 U4506 ( .A1(n3774), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[22][26] ), .B2(n3773), .ZN(n4874) );
  OAI22_X1 U4507 ( .A1(n3774), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[22][27] ), .B2(n3772), .ZN(n4875) );
  OAI22_X1 U4508 ( .A1(n3774), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[22][28] ), .B2(n3773), .ZN(n4876) );
  OAI22_X1 U4509 ( .A1(n3774), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[22][29] ), .B2(n3772), .ZN(n4877) );
  OAI22_X1 U4510 ( .A1(n3774), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[22][30] ), .B2(n3773), .ZN(n4878) );
  OAI22_X1 U4511 ( .A1(n3774), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[22][31] ), .B2(n3773), .ZN(n4879) );
  NOR2_X2 U4512 ( .A1(n3891), .A2(n3775), .ZN(n3776) );
  INV_X2 U4513 ( .A(n3777), .ZN(n3778) );
  OAI22_X1 U4514 ( .A1(n3778), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[23][0] ), .B2(n3777), .ZN(n4880) );
  OAI22_X1 U4515 ( .A1(n3778), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[23][1] ), .B2(n3776), .ZN(n4881) );
  OAI22_X1 U4516 ( .A1(n3778), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[23][2] ), .B2(n3776), .ZN(n4882) );
  OAI22_X1 U4517 ( .A1(n3778), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[23][3] ), .B2(n3776), .ZN(n4883) );
  OAI22_X1 U4518 ( .A1(n3778), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[23][4] ), .B2(n3776), .ZN(n4884) );
  OAI22_X1 U4519 ( .A1(n3778), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[23][5] ), .B2(n3776), .ZN(n4885) );
  OAI22_X1 U4520 ( .A1(n3778), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[23][6] ), .B2(n3776), .ZN(n4886) );
  OAI22_X1 U4521 ( .A1(n3778), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[23][7] ), .B2(n3776), .ZN(n4887) );
  OAI22_X1 U4522 ( .A1(n3778), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[23][8] ), .B2(n3776), .ZN(n4888) );
  OAI22_X1 U4523 ( .A1(n3778), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[23][9] ), .B2(n3776), .ZN(n4889) );
  OAI22_X1 U4524 ( .A1(n3778), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[23][10] ), .B2(n3776), .ZN(n4890) );
  OAI22_X1 U4525 ( .A1(n3778), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[23][11] ), .B2(n3776), .ZN(n4891) );
  OAI22_X1 U4526 ( .A1(n3778), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[23][12] ), .B2(n3776), .ZN(n4892) );
  OAI22_X1 U4527 ( .A1(n3778), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[23][13] ), .B2(n3776), .ZN(n4893) );
  OAI22_X1 U4528 ( .A1(n3778), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[23][14] ), .B2(n3776), .ZN(n4894) );
  OAI22_X1 U4529 ( .A1(n3778), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[23][15] ), .B2(n3777), .ZN(n4895) );
  OAI22_X1 U4530 ( .A1(n3778), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[23][16] ), .B2(n3776), .ZN(n4896) );
  OAI22_X1 U4531 ( .A1(n3778), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[23][17] ), .B2(n3776), .ZN(n4897) );
  OAI22_X1 U4532 ( .A1(n3778), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[23][18] ), .B2(n3776), .ZN(n4898) );
  OAI22_X1 U4533 ( .A1(n3778), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[23][19] ), .B2(n3777), .ZN(n4899) );
  OAI22_X1 U4534 ( .A1(n3778), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[23][20] ), .B2(n3776), .ZN(n4900) );
  OAI22_X1 U4535 ( .A1(n3778), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[23][21] ), .B2(n3776), .ZN(n4901) );
  OAI22_X1 U4536 ( .A1(n3778), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[23][22] ), .B2(n3777), .ZN(n4902) );
  OAI22_X1 U4537 ( .A1(n3778), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[23][23] ), .B2(n3777), .ZN(n4903) );
  OAI22_X1 U4538 ( .A1(n3778), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[23][24] ), .B2(n3777), .ZN(n4904) );
  OAI22_X1 U4539 ( .A1(n3778), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[23][25] ), .B2(n3776), .ZN(n4905) );
  OAI22_X1 U4540 ( .A1(n3778), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[23][26] ), .B2(n3777), .ZN(n4906) );
  OAI22_X1 U4541 ( .A1(n3778), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[23][27] ), .B2(n3776), .ZN(n4907) );
  OAI22_X1 U4542 ( .A1(n3778), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[23][28] ), .B2(n3777), .ZN(n4908) );
  OAI22_X1 U4543 ( .A1(n3778), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[23][29] ), .B2(n3776), .ZN(n4909) );
  OAI22_X1 U4544 ( .A1(n3778), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[23][30] ), .B2(n3777), .ZN(n4910) );
  OAI22_X1 U4545 ( .A1(n3778), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[23][31] ), .B2(n3777), .ZN(n4911) );
  NOR2_X2 U4546 ( .A1(n3897), .A2(n3801), .ZN(n3780) );
  INV_X2 U4547 ( .A(n3781), .ZN(n3782) );
  OAI22_X1 U4548 ( .A1(n3782), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[24][0] ), .B2(n3781), .ZN(n4912) );
  OAI22_X1 U4549 ( .A1(n3782), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[24][1] ), .B2(n3780), .ZN(n4913) );
  OAI22_X1 U4550 ( .A1(n3782), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[24][2] ), .B2(n3780), .ZN(n4914) );
  OAI22_X1 U4551 ( .A1(n3782), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[24][3] ), .B2(n3780), .ZN(n4915) );
  OAI22_X1 U4552 ( .A1(n3782), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[24][4] ), .B2(n3780), .ZN(n4916) );
  OAI22_X1 U4553 ( .A1(n3782), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[24][5] ), .B2(n3780), .ZN(n4917) );
  OAI22_X1 U4554 ( .A1(n3782), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[24][6] ), .B2(n3780), .ZN(n4918) );
  OAI22_X1 U4555 ( .A1(n3782), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[24][7] ), .B2(n3780), .ZN(n4919) );
  OAI22_X1 U4556 ( .A1(n3782), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[24][8] ), .B2(n3780), .ZN(n4920) );
  OAI22_X1 U4557 ( .A1(n3782), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[24][9] ), .B2(n3780), .ZN(n4921) );
  OAI22_X1 U4558 ( .A1(n3782), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[24][10] ), .B2(n3780), .ZN(n4922) );
  OAI22_X1 U4559 ( .A1(n3782), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[24][11] ), .B2(n3780), .ZN(n4923) );
  OAI22_X1 U4560 ( .A1(n3782), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[24][12] ), .B2(n3780), .ZN(n4924) );
  OAI22_X1 U4561 ( .A1(n3782), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[24][13] ), .B2(n3780), .ZN(n4925) );
  OAI22_X1 U4562 ( .A1(n3782), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[24][14] ), .B2(n3780), .ZN(n4926) );
  OAI22_X1 U4563 ( .A1(n3782), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[24][15] ), .B2(n3781), .ZN(n4927) );
  OAI22_X1 U4564 ( .A1(n3782), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[24][16] ), .B2(n3780), .ZN(n4928) );
  OAI22_X1 U4565 ( .A1(n3782), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[24][17] ), .B2(n3780), .ZN(n4929) );
  OAI22_X1 U4566 ( .A1(n3782), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[24][18] ), .B2(n3780), .ZN(n4930) );
  OAI22_X1 U4567 ( .A1(n3782), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[24][19] ), .B2(n3781), .ZN(n4931) );
  OAI22_X1 U4568 ( .A1(n3782), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[24][20] ), .B2(n3780), .ZN(n4932) );
  OAI22_X1 U4569 ( .A1(n3782), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[24][21] ), .B2(n3780), .ZN(n4933) );
  OAI22_X1 U4570 ( .A1(n3782), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[24][22] ), .B2(n3781), .ZN(n4934) );
  OAI22_X1 U4571 ( .A1(n3782), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[24][23] ), .B2(n3781), .ZN(n4935) );
  OAI22_X1 U4572 ( .A1(n3782), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[24][24] ), .B2(n3781), .ZN(n4936) );
  OAI22_X1 U4573 ( .A1(n3782), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[24][25] ), .B2(n3780), .ZN(n4937) );
  OAI22_X1 U4574 ( .A1(n3782), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[24][26] ), .B2(n3781), .ZN(n4938) );
  OAI22_X1 U4575 ( .A1(n3782), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[24][27] ), .B2(n3780), .ZN(n4939) );
  OAI22_X1 U4576 ( .A1(n3782), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[24][28] ), .B2(n3781), .ZN(n4940) );
  OAI22_X1 U4577 ( .A1(n3782), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[24][29] ), .B2(n3780), .ZN(n4941) );
  OAI22_X1 U4578 ( .A1(n3782), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[24][30] ), .B2(n3781), .ZN(n4942) );
  OAI22_X1 U4579 ( .A1(n3782), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[24][31] ), .B2(n3781), .ZN(n4943) );
  NOR2_X2 U4580 ( .A1(n3933), .A2(n3801), .ZN(n3783) );
  INV_X2 U4581 ( .A(n3784), .ZN(n3785) );
  OAI22_X1 U4582 ( .A1(n3785), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[25][0] ), .B2(n3784), .ZN(n4944) );
  OAI22_X1 U4583 ( .A1(n3785), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[25][1] ), .B2(n3783), .ZN(n4945) );
  OAI22_X1 U4584 ( .A1(n3785), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[25][2] ), .B2(n3783), .ZN(n4946) );
  OAI22_X1 U4585 ( .A1(n3785), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[25][3] ), .B2(n3783), .ZN(n4947) );
  OAI22_X1 U4586 ( .A1(n3785), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[25][4] ), .B2(n3783), .ZN(n4948) );
  OAI22_X1 U4587 ( .A1(n3785), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[25][5] ), .B2(n3783), .ZN(n4949) );
  OAI22_X1 U4588 ( .A1(n3785), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[25][6] ), .B2(n3783), .ZN(n4950) );
  OAI22_X1 U4589 ( .A1(n3785), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[25][7] ), .B2(n3783), .ZN(n4951) );
  OAI22_X1 U4590 ( .A1(n3785), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[25][8] ), .B2(n3783), .ZN(n4952) );
  OAI22_X1 U4591 ( .A1(n3785), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[25][9] ), .B2(n3783), .ZN(n4953) );
  OAI22_X1 U4592 ( .A1(n3785), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[25][10] ), .B2(n3783), .ZN(n4954) );
  OAI22_X1 U4593 ( .A1(n3785), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[25][11] ), .B2(n3783), .ZN(n4955) );
  OAI22_X1 U4594 ( .A1(n3785), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[25][12] ), .B2(n3783), .ZN(n4956) );
  OAI22_X1 U4595 ( .A1(n3785), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[25][13] ), .B2(n3783), .ZN(n4957) );
  OAI22_X1 U4596 ( .A1(n3785), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[25][14] ), .B2(n3783), .ZN(n4958) );
  OAI22_X1 U4597 ( .A1(n3785), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[25][15] ), .B2(n3784), .ZN(n4959) );
  OAI22_X1 U4598 ( .A1(n3785), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[25][16] ), .B2(n3783), .ZN(n4960) );
  OAI22_X1 U4599 ( .A1(n3785), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[25][17] ), .B2(n3783), .ZN(n4961) );
  OAI22_X1 U4600 ( .A1(n3785), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[25][18] ), .B2(n3783), .ZN(n4962) );
  OAI22_X1 U4601 ( .A1(n3785), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[25][19] ), .B2(n3784), .ZN(n4963) );
  OAI22_X1 U4602 ( .A1(n3785), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[25][20] ), .B2(n3783), .ZN(n4964) );
  OAI22_X1 U4603 ( .A1(n3785), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[25][21] ), .B2(n3783), .ZN(n4965) );
  OAI22_X1 U4604 ( .A1(n3785), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[25][22] ), .B2(n3784), .ZN(n4966) );
  OAI22_X1 U4605 ( .A1(n3785), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[25][23] ), .B2(n3784), .ZN(n4967) );
  OAI22_X1 U4606 ( .A1(n3785), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[25][24] ), .B2(n3784), .ZN(n4968) );
  OAI22_X1 U4607 ( .A1(n3785), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[25][25] ), .B2(n3783), .ZN(n4969) );
  OAI22_X1 U4608 ( .A1(n3785), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[25][26] ), .B2(n3784), .ZN(n4970) );
  OAI22_X1 U4609 ( .A1(n3785), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[25][27] ), .B2(n3783), .ZN(n4971) );
  OAI22_X1 U4610 ( .A1(n3785), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[25][28] ), .B2(n3784), .ZN(n4972) );
  OAI22_X1 U4611 ( .A1(n3785), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[25][29] ), .B2(n3783), .ZN(n4973) );
  OAI22_X1 U4612 ( .A1(n3785), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[25][30] ), .B2(n3784), .ZN(n4974) );
  OAI22_X1 U4613 ( .A1(n3785), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[25][31] ), .B2(n3784), .ZN(n4975) );
  NOR2_X2 U4614 ( .A1(n3970), .A2(n3801), .ZN(n3786) );
  INV_X2 U4615 ( .A(n3787), .ZN(n3788) );
  OAI22_X1 U4616 ( .A1(n3788), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[26][0] ), .B2(n3787), .ZN(n4976) );
  OAI22_X1 U4617 ( .A1(n3788), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[26][1] ), .B2(n3786), .ZN(n4977) );
  OAI22_X1 U4618 ( .A1(n3788), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[26][2] ), .B2(n3786), .ZN(n4978) );
  OAI22_X1 U4619 ( .A1(n3788), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[26][3] ), .B2(n3786), .ZN(n4979) );
  OAI22_X1 U4620 ( .A1(n3788), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[26][4] ), .B2(n3786), .ZN(n4980) );
  OAI22_X1 U4621 ( .A1(n3788), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[26][5] ), .B2(n3786), .ZN(n4981) );
  OAI22_X1 U4622 ( .A1(n3788), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[26][6] ), .B2(n3786), .ZN(n4982) );
  OAI22_X1 U4623 ( .A1(n3788), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[26][7] ), .B2(n3786), .ZN(n4983) );
  OAI22_X1 U4624 ( .A1(n3788), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[26][8] ), .B2(n3786), .ZN(n4984) );
  OAI22_X1 U4625 ( .A1(n3788), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[26][9] ), .B2(n3786), .ZN(n4985) );
  OAI22_X1 U4626 ( .A1(n3788), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[26][10] ), .B2(n3786), .ZN(n4986) );
  OAI22_X1 U4627 ( .A1(n3788), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[26][11] ), .B2(n3786), .ZN(n4987) );
  OAI22_X1 U4628 ( .A1(n3788), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[26][12] ), .B2(n3786), .ZN(n4988) );
  OAI22_X1 U4629 ( .A1(n3788), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[26][13] ), .B2(n3786), .ZN(n4989) );
  OAI22_X1 U4630 ( .A1(n3788), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[26][14] ), .B2(n3786), .ZN(n4990) );
  OAI22_X1 U4631 ( .A1(n3788), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[26][15] ), .B2(n3787), .ZN(n4991) );
  OAI22_X1 U4632 ( .A1(n3788), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[26][16] ), .B2(n3786), .ZN(n4992) );
  OAI22_X1 U4633 ( .A1(n3788), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[26][17] ), .B2(n3786), .ZN(n4993) );
  OAI22_X1 U4634 ( .A1(n3788), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[26][18] ), .B2(n3786), .ZN(n4994) );
  OAI22_X1 U4635 ( .A1(n3788), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[26][19] ), .B2(n3787), .ZN(n4995) );
  OAI22_X1 U4636 ( .A1(n3788), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[26][20] ), .B2(n3786), .ZN(n4996) );
  OAI22_X1 U4637 ( .A1(n3788), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[26][21] ), .B2(n3786), .ZN(n4997) );
  OAI22_X1 U4638 ( .A1(n3788), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[26][22] ), .B2(n3787), .ZN(n4998) );
  OAI22_X1 U4639 ( .A1(n3788), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[26][23] ), .B2(n3787), .ZN(n4999) );
  OAI22_X1 U4640 ( .A1(n3788), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[26][24] ), .B2(n3787), .ZN(n5000) );
  OAI22_X1 U4641 ( .A1(n3788), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[26][25] ), .B2(n3786), .ZN(n5001) );
  OAI22_X1 U4642 ( .A1(n3788), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[26][26] ), .B2(n3787), .ZN(n5002) );
  OAI22_X1 U4643 ( .A1(n3788), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[26][27] ), .B2(n3786), .ZN(n5003) );
  OAI22_X1 U4644 ( .A1(n3788), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[26][28] ), .B2(n3787), .ZN(n5004) );
  OAI22_X1 U4645 ( .A1(n3788), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[26][29] ), .B2(n3786), .ZN(n5005) );
  OAI22_X1 U4646 ( .A1(n3788), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[26][30] ), .B2(n3787), .ZN(n5006) );
  OAI22_X1 U4647 ( .A1(n3788), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[26][31] ), .B2(n3787), .ZN(n5007) );
  NOR2_X2 U4648 ( .A1(n3873), .A2(n3801), .ZN(n3789) );
  INV_X2 U4649 ( .A(n3790), .ZN(n3791) );
  OAI22_X1 U4650 ( .A1(n3791), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[27][0] ), .B2(n3790), .ZN(n5008) );
  OAI22_X1 U4651 ( .A1(n3791), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[27][1] ), .B2(n3789), .ZN(n5009) );
  OAI22_X1 U4652 ( .A1(n3791), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[27][2] ), .B2(n3789), .ZN(n5010) );
  OAI22_X1 U4653 ( .A1(n3791), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[27][3] ), .B2(n3789), .ZN(n5011) );
  OAI22_X1 U4654 ( .A1(n3791), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[27][4] ), .B2(n3789), .ZN(n5012) );
  OAI22_X1 U4655 ( .A1(n3791), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[27][5] ), .B2(n3789), .ZN(n5013) );
  OAI22_X1 U4656 ( .A1(n3791), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[27][6] ), .B2(n3789), .ZN(n5014) );
  OAI22_X1 U4657 ( .A1(n3791), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[27][7] ), .B2(n3789), .ZN(n5015) );
  OAI22_X1 U4658 ( .A1(n3791), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[27][8] ), .B2(n3789), .ZN(n5016) );
  OAI22_X1 U4659 ( .A1(n3791), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[27][9] ), .B2(n3789), .ZN(n5017) );
  OAI22_X1 U4660 ( .A1(n3791), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[27][10] ), .B2(n3789), .ZN(n5018) );
  OAI22_X1 U4661 ( .A1(n3791), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[27][11] ), .B2(n3789), .ZN(n5019) );
  OAI22_X1 U4662 ( .A1(n3791), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[27][12] ), .B2(n3789), .ZN(n5020) );
  OAI22_X1 U4663 ( .A1(n3791), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[27][13] ), .B2(n3789), .ZN(n5021) );
  OAI22_X1 U4664 ( .A1(n3791), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[27][14] ), .B2(n3789), .ZN(n5022) );
  OAI22_X1 U4665 ( .A1(n3791), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[27][15] ), .B2(n3790), .ZN(n5023) );
  OAI22_X1 U4666 ( .A1(n3791), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[27][16] ), .B2(n3789), .ZN(n5024) );
  OAI22_X1 U4667 ( .A1(n3791), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[27][17] ), .B2(n3789), .ZN(n5025) );
  OAI22_X1 U4668 ( .A1(n3791), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[27][18] ), .B2(n3789), .ZN(n5026) );
  OAI22_X1 U4669 ( .A1(n3791), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[27][19] ), .B2(n3790), .ZN(n5027) );
  OAI22_X1 U4670 ( .A1(n3791), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[27][20] ), .B2(n3789), .ZN(n5028) );
  OAI22_X1 U4671 ( .A1(n3791), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[27][21] ), .B2(n3789), .ZN(n5029) );
  OAI22_X1 U4672 ( .A1(n3791), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[27][22] ), .B2(n3790), .ZN(n5030) );
  OAI22_X1 U4673 ( .A1(n3791), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[27][23] ), .B2(n3790), .ZN(n5031) );
  OAI22_X1 U4674 ( .A1(n3791), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[27][24] ), .B2(n3790), .ZN(n5032) );
  OAI22_X1 U4675 ( .A1(n3791), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[27][25] ), .B2(n3789), .ZN(n5033) );
  OAI22_X1 U4676 ( .A1(n3791), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[27][26] ), .B2(n3790), .ZN(n5034) );
  OAI22_X1 U4677 ( .A1(n3791), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[27][27] ), .B2(n3789), .ZN(n5035) );
  OAI22_X1 U4678 ( .A1(n3791), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[27][28] ), .B2(n3790), .ZN(n5036) );
  OAI22_X1 U4679 ( .A1(n3791), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[27][29] ), .B2(n3789), .ZN(n5037) );
  OAI22_X1 U4680 ( .A1(n3791), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[27][30] ), .B2(n3790), .ZN(n5038) );
  OAI22_X1 U4681 ( .A1(n3791), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[27][31] ), .B2(n3790), .ZN(n5039) );
  NOR2_X2 U4682 ( .A1(n3878), .A2(n3801), .ZN(n3792) );
  INV_X2 U4683 ( .A(n3793), .ZN(n3794) );
  OAI22_X1 U4684 ( .A1(n3794), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[28][0] ), .B2(n3793), .ZN(n5040) );
  OAI22_X1 U4685 ( .A1(n3794), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[28][1] ), .B2(n3792), .ZN(n5041) );
  OAI22_X1 U4686 ( .A1(n3794), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[28][2] ), .B2(n3792), .ZN(n5042) );
  OAI22_X1 U4687 ( .A1(n3794), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[28][3] ), .B2(n3792), .ZN(n5043) );
  OAI22_X1 U4688 ( .A1(n3794), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[28][4] ), .B2(n3792), .ZN(n5044) );
  OAI22_X1 U4689 ( .A1(n3794), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[28][5] ), .B2(n3792), .ZN(n5045) );
  OAI22_X1 U4690 ( .A1(n3794), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[28][6] ), .B2(n3792), .ZN(n5046) );
  OAI22_X1 U4691 ( .A1(n3794), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[28][7] ), .B2(n3792), .ZN(n5047) );
  OAI22_X1 U4692 ( .A1(n3794), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[28][8] ), .B2(n3792), .ZN(n5048) );
  OAI22_X1 U4693 ( .A1(n3794), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[28][9] ), .B2(n3792), .ZN(n5049) );
  OAI22_X1 U4694 ( .A1(n3794), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[28][10] ), .B2(n3792), .ZN(n5050) );
  OAI22_X1 U4695 ( .A1(n3794), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[28][11] ), .B2(n3792), .ZN(n5051) );
  OAI22_X1 U4696 ( .A1(n3794), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[28][12] ), .B2(n3792), .ZN(n5052) );
  OAI22_X1 U4697 ( .A1(n3794), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[28][13] ), .B2(n3792), .ZN(n5053) );
  OAI22_X1 U4698 ( .A1(n3794), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[28][14] ), .B2(n3792), .ZN(n5054) );
  OAI22_X1 U4699 ( .A1(n3794), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[28][15] ), .B2(n3793), .ZN(n5055) );
  OAI22_X1 U4700 ( .A1(n3794), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[28][16] ), .B2(n3792), .ZN(n5056) );
  OAI22_X1 U4701 ( .A1(n3794), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[28][17] ), .B2(n3792), .ZN(n5057) );
  OAI22_X1 U4702 ( .A1(n3794), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[28][18] ), .B2(n3792), .ZN(n5058) );
  OAI22_X1 U4703 ( .A1(n3794), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[28][19] ), .B2(n3793), .ZN(n5059) );
  OAI22_X1 U4704 ( .A1(n3794), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[28][20] ), .B2(n3792), .ZN(n5060) );
  OAI22_X1 U4705 ( .A1(n3794), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[28][21] ), .B2(n3792), .ZN(n5061) );
  OAI22_X1 U4706 ( .A1(n3794), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[28][22] ), .B2(n3793), .ZN(n5062) );
  OAI22_X1 U4707 ( .A1(n3794), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[28][23] ), .B2(n3793), .ZN(n5063) );
  OAI22_X1 U4708 ( .A1(n3794), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[28][24] ), .B2(n3793), .ZN(n5064) );
  OAI22_X1 U4709 ( .A1(n3794), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[28][25] ), .B2(n3792), .ZN(n5065) );
  OAI22_X1 U4710 ( .A1(n3794), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[28][26] ), .B2(n3793), .ZN(n5066) );
  OAI22_X1 U4711 ( .A1(n3794), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[28][27] ), .B2(n3792), .ZN(n5067) );
  OAI22_X1 U4712 ( .A1(n3794), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[28][28] ), .B2(n3793), .ZN(n5068) );
  OAI22_X1 U4713 ( .A1(n3794), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[28][29] ), .B2(n3792), .ZN(n5069) );
  OAI22_X1 U4714 ( .A1(n3794), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[28][30] ), .B2(n3793), .ZN(n5070) );
  OAI22_X1 U4715 ( .A1(n3794), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[28][31] ), .B2(n3793), .ZN(n5071) );
  NOR2_X2 U4716 ( .A1(n3882), .A2(n3801), .ZN(n3795) );
  INV_X2 U4717 ( .A(n3796), .ZN(n3797) );
  OAI22_X1 U4718 ( .A1(n3797), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[29][0] ), .B2(n3796), .ZN(n5072) );
  OAI22_X1 U4719 ( .A1(n3797), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[29][1] ), .B2(n3795), .ZN(n5073) );
  OAI22_X1 U4720 ( .A1(n3797), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[29][2] ), .B2(n3795), .ZN(n5074) );
  OAI22_X1 U4721 ( .A1(n3797), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[29][3] ), .B2(n3795), .ZN(n5075) );
  OAI22_X1 U4722 ( .A1(n3797), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[29][4] ), .B2(n3795), .ZN(n5076) );
  OAI22_X1 U4723 ( .A1(n3797), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[29][5] ), .B2(n3795), .ZN(n5077) );
  OAI22_X1 U4724 ( .A1(n3797), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[29][6] ), .B2(n3795), .ZN(n5078) );
  OAI22_X1 U4725 ( .A1(n3797), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[29][7] ), .B2(n3795), .ZN(n5079) );
  OAI22_X1 U4726 ( .A1(n3797), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[29][8] ), .B2(n3795), .ZN(n5080) );
  OAI22_X1 U4727 ( .A1(n3797), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[29][9] ), .B2(n3795), .ZN(n5081) );
  OAI22_X1 U4728 ( .A1(n3797), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[29][10] ), .B2(n3795), .ZN(n5082) );
  OAI22_X1 U4729 ( .A1(n3797), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[29][11] ), .B2(n3795), .ZN(n5083) );
  OAI22_X1 U4730 ( .A1(n3797), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[29][12] ), .B2(n3795), .ZN(n5084) );
  OAI22_X1 U4731 ( .A1(n3797), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[29][13] ), .B2(n3795), .ZN(n5085) );
  OAI22_X1 U4732 ( .A1(n3797), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[29][14] ), .B2(n3795), .ZN(n5086) );
  OAI22_X1 U4733 ( .A1(n3797), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[29][15] ), .B2(n3796), .ZN(n5087) );
  OAI22_X1 U4734 ( .A1(n3797), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[29][16] ), .B2(n3795), .ZN(n5088) );
  OAI22_X1 U4735 ( .A1(n3797), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[29][17] ), .B2(n3795), .ZN(n5089) );
  OAI22_X1 U4736 ( .A1(n3797), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[29][18] ), .B2(n3795), .ZN(n5090) );
  OAI22_X1 U4737 ( .A1(n3797), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[29][19] ), .B2(n3796), .ZN(n5091) );
  OAI22_X1 U4738 ( .A1(n3797), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[29][20] ), .B2(n3795), .ZN(n5092) );
  OAI22_X1 U4739 ( .A1(n3797), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[29][21] ), .B2(n3795), .ZN(n5093) );
  OAI22_X1 U4740 ( .A1(n3797), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[29][22] ), .B2(n3796), .ZN(n5094) );
  OAI22_X1 U4741 ( .A1(n3797), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[29][23] ), .B2(n3796), .ZN(n5095) );
  OAI22_X1 U4742 ( .A1(n3797), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[29][24] ), .B2(n3796), .ZN(n5096) );
  OAI22_X1 U4743 ( .A1(n3797), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[29][25] ), .B2(n3795), .ZN(n5097) );
  OAI22_X1 U4744 ( .A1(n3797), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[29][26] ), .B2(n3796), .ZN(n5098) );
  OAI22_X1 U4745 ( .A1(n3797), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[29][27] ), .B2(n3795), .ZN(n5099) );
  OAI22_X1 U4746 ( .A1(n3797), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[29][28] ), .B2(n3796), .ZN(n5100) );
  OAI22_X1 U4747 ( .A1(n3797), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[29][29] ), .B2(n3795), .ZN(n5101) );
  OAI22_X1 U4748 ( .A1(n3797), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[29][30] ), .B2(n3796), .ZN(n5102) );
  OAI22_X1 U4749 ( .A1(n3797), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[29][31] ), .B2(n3796), .ZN(n5103) );
  NOR2_X2 U4750 ( .A1(n3886), .A2(n3801), .ZN(n3798) );
  INV_X2 U4751 ( .A(n3799), .ZN(n3800) );
  OAI22_X1 U4752 ( .A1(n3800), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[30][0] ), .B2(n3799), .ZN(n5104) );
  OAI22_X1 U4753 ( .A1(n3800), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[30][1] ), .B2(n3798), .ZN(n5105) );
  OAI22_X1 U4754 ( .A1(n3800), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[30][2] ), .B2(n3798), .ZN(n5106) );
  OAI22_X1 U4755 ( .A1(n3800), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[30][3] ), .B2(n3798), .ZN(n5107) );
  OAI22_X1 U4756 ( .A1(n3800), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[30][4] ), .B2(n3798), .ZN(n5108) );
  OAI22_X1 U4757 ( .A1(n3800), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[30][5] ), .B2(n3798), .ZN(n5109) );
  OAI22_X1 U4758 ( .A1(n3800), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[30][6] ), .B2(n3798), .ZN(n5110) );
  OAI22_X1 U4759 ( .A1(n3800), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[30][7] ), .B2(n3798), .ZN(n5111) );
  OAI22_X1 U4760 ( .A1(n3800), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[30][8] ), .B2(n3798), .ZN(n5112) );
  OAI22_X1 U4761 ( .A1(n3800), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[30][9] ), .B2(n3798), .ZN(n5113) );
  OAI22_X1 U4762 ( .A1(n3800), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[30][10] ), .B2(n3798), .ZN(n5114) );
  OAI22_X1 U4763 ( .A1(n3800), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[30][11] ), .B2(n3798), .ZN(n5115) );
  OAI22_X1 U4764 ( .A1(n3800), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[30][12] ), .B2(n3798), .ZN(n5116) );
  OAI22_X1 U4765 ( .A1(n3800), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[30][13] ), .B2(n3798), .ZN(n5117) );
  OAI22_X1 U4766 ( .A1(n3800), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[30][14] ), .B2(n3798), .ZN(n5118) );
  OAI22_X1 U4767 ( .A1(n3800), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[30][15] ), .B2(n3799), .ZN(n5119) );
  OAI22_X1 U4768 ( .A1(n3800), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[30][16] ), .B2(n3798), .ZN(n5120) );
  OAI22_X1 U4769 ( .A1(n3800), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[30][17] ), .B2(n3798), .ZN(n5121) );
  OAI22_X1 U4770 ( .A1(n3800), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[30][18] ), .B2(n3798), .ZN(n5122) );
  OAI22_X1 U4771 ( .A1(n3800), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[30][19] ), .B2(n3799), .ZN(n5123) );
  OAI22_X1 U4772 ( .A1(n3800), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[30][20] ), .B2(n3798), .ZN(n5124) );
  OAI22_X1 U4773 ( .A1(n3800), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[30][21] ), .B2(n3798), .ZN(n5125) );
  OAI22_X1 U4774 ( .A1(n3800), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[30][22] ), .B2(n3799), .ZN(n5126) );
  OAI22_X1 U4775 ( .A1(n3800), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[30][23] ), .B2(n3799), .ZN(n5127) );
  OAI22_X1 U4776 ( .A1(n3800), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[30][24] ), .B2(n3799), .ZN(n5128) );
  OAI22_X1 U4777 ( .A1(n3800), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[30][25] ), .B2(n3798), .ZN(n5129) );
  OAI22_X1 U4778 ( .A1(n3800), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[30][26] ), .B2(n3799), .ZN(n5130) );
  OAI22_X1 U4779 ( .A1(n3800), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[30][27] ), .B2(n3798), .ZN(n5131) );
  OAI22_X1 U4780 ( .A1(n3800), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[30][28] ), .B2(n3799), .ZN(n5132) );
  OAI22_X1 U4781 ( .A1(n3800), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[30][29] ), .B2(n3798), .ZN(n5133) );
  OAI22_X1 U4782 ( .A1(n3800), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[30][30] ), .B2(n3799), .ZN(n5134) );
  OAI22_X1 U4783 ( .A1(n3800), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[30][31] ), .B2(n3799), .ZN(n5135) );
  NOR2_X2 U4784 ( .A1(n3891), .A2(n3801), .ZN(n3802) );
  INV_X2 U4785 ( .A(n3803), .ZN(n3804) );
  OAI22_X1 U4786 ( .A1(n3804), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[31][0] ), .B2(n3803), .ZN(n5136) );
  OAI22_X1 U4787 ( .A1(n3804), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[31][1] ), .B2(n3802), .ZN(n5137) );
  OAI22_X1 U4788 ( .A1(n3804), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[31][2] ), .B2(n3802), .ZN(n5138) );
  OAI22_X1 U4789 ( .A1(n3804), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[31][3] ), .B2(n3802), .ZN(n5139) );
  OAI22_X1 U4790 ( .A1(n3804), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[31][4] ), .B2(n3802), .ZN(n5140) );
  OAI22_X1 U4791 ( .A1(n3804), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[31][5] ), .B2(n3802), .ZN(n5141) );
  OAI22_X1 U4792 ( .A1(n3804), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[31][6] ), .B2(n3802), .ZN(n5142) );
  OAI22_X1 U4793 ( .A1(n3804), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[31][7] ), .B2(n3802), .ZN(n5143) );
  OAI22_X1 U4794 ( .A1(n3804), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[31][8] ), .B2(n3802), .ZN(n5144) );
  OAI22_X1 U4795 ( .A1(n3804), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[31][9] ), .B2(n3802), .ZN(n5145) );
  OAI22_X1 U4796 ( .A1(n3804), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[31][10] ), .B2(n3802), .ZN(n5146) );
  OAI22_X1 U4797 ( .A1(n3804), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[31][11] ), .B2(n3802), .ZN(n5147) );
  OAI22_X1 U4798 ( .A1(n3804), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[31][12] ), .B2(n3802), .ZN(n5148) );
  OAI22_X1 U4799 ( .A1(n3804), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[31][13] ), .B2(n3802), .ZN(n5149) );
  OAI22_X1 U4800 ( .A1(n3804), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[31][14] ), .B2(n3802), .ZN(n5150) );
  OAI22_X1 U4801 ( .A1(n3804), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[31][15] ), .B2(n3803), .ZN(n5151) );
  OAI22_X1 U4802 ( .A1(n3804), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[31][16] ), .B2(n3802), .ZN(n5152) );
  OAI22_X1 U4803 ( .A1(n3804), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[31][17] ), .B2(n3802), .ZN(n5153) );
  OAI22_X1 U4804 ( .A1(n3804), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[31][18] ), .B2(n3802), .ZN(n5154) );
  OAI22_X1 U4805 ( .A1(n3804), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[31][19] ), .B2(n3803), .ZN(n5155) );
  OAI22_X1 U4806 ( .A1(n3804), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[31][20] ), .B2(n3802), .ZN(n5156) );
  OAI22_X1 U4807 ( .A1(n3804), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[31][21] ), .B2(n3802), .ZN(n5157) );
  OAI22_X1 U4808 ( .A1(n3804), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[31][22] ), .B2(n3803), .ZN(n5158) );
  OAI22_X1 U4809 ( .A1(n3804), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[31][23] ), .B2(n3803), .ZN(n5159) );
  OAI22_X1 U4810 ( .A1(n3804), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[31][24] ), .B2(n3803), .ZN(n5160) );
  OAI22_X1 U4811 ( .A1(n3804), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[31][25] ), .B2(n3802), .ZN(n5161) );
  OAI22_X1 U4812 ( .A1(n3804), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[31][26] ), .B2(n3803), .ZN(n5162) );
  OAI22_X1 U4813 ( .A1(n3804), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[31][27] ), .B2(n3802), .ZN(n5163) );
  OAI22_X1 U4814 ( .A1(n3804), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[31][28] ), .B2(n3803), .ZN(n5164) );
  OAI22_X1 U4815 ( .A1(n3804), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[31][29] ), .B2(n3802), .ZN(n5165) );
  OAI22_X1 U4816 ( .A1(n3804), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[31][30] ), .B2(n3803), .ZN(n5166) );
  OAI22_X1 U4817 ( .A1(n3804), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[31][31] ), .B2(n3803), .ZN(n5167) );
  NOR2_X2 U4818 ( .A1(n3897), .A2(n3890), .ZN(n3832) );
  INV_X2 U4819 ( .A(n3834), .ZN(n3835) );
  OAI22_X1 U4820 ( .A1(n3835), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[32][0] ), .B2(n3834), .ZN(n3805) );
  INV_X1 U4821 ( .A(n3805), .ZN(\xmem_inst/n3466 ) );
  OAI22_X1 U4822 ( .A1(n3835), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[32][1] ), .B2(n3832), .ZN(n3806) );
  INV_X1 U4823 ( .A(n3806), .ZN(\xmem_inst/n3467 ) );
  OAI22_X1 U4824 ( .A1(n3835), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[32][2] ), .B2(n3832), .ZN(n3807) );
  INV_X1 U4825 ( .A(n3807), .ZN(\xmem_inst/n3468 ) );
  OAI22_X1 U4826 ( .A1(n3835), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[32][3] ), .B2(n3832), .ZN(n3808) );
  INV_X1 U4827 ( .A(n3808), .ZN(\xmem_inst/n3469 ) );
  OAI22_X1 U4828 ( .A1(n3835), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[32][4] ), .B2(n3832), .ZN(n3809) );
  INV_X1 U4829 ( .A(n3809), .ZN(\xmem_inst/n3470 ) );
  OAI22_X1 U4830 ( .A1(n3835), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[32][5] ), .B2(n3832), .ZN(n3810) );
  INV_X1 U4831 ( .A(n3810), .ZN(\xmem_inst/n3471 ) );
  OAI22_X1 U4832 ( .A1(n3835), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[32][6] ), .B2(n3832), .ZN(n3811) );
  INV_X1 U4833 ( .A(n3811), .ZN(\xmem_inst/n3472 ) );
  OAI22_X1 U4834 ( .A1(n3835), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[32][7] ), .B2(n3832), .ZN(n3812) );
  INV_X1 U4835 ( .A(n3812), .ZN(\xmem_inst/n3473 ) );
  OAI22_X1 U4836 ( .A1(n3835), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[32][8] ), .B2(n3832), .ZN(n3813) );
  INV_X1 U4837 ( .A(n3813), .ZN(\xmem_inst/n3474 ) );
  OAI22_X1 U4838 ( .A1(n3835), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[32][9] ), .B2(n3832), .ZN(n3814) );
  INV_X1 U4839 ( .A(n3814), .ZN(\xmem_inst/n3475 ) );
  OAI22_X1 U4840 ( .A1(n3835), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[32][10] ), .B2(n3832), .ZN(n3815) );
  INV_X1 U4841 ( .A(n3815), .ZN(\xmem_inst/n3476 ) );
  OAI22_X1 U4842 ( .A1(n3835), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[32][11] ), .B2(n3832), .ZN(n3816) );
  INV_X1 U4843 ( .A(n3816), .ZN(\xmem_inst/n3477 ) );
  OAI22_X1 U4844 ( .A1(n3835), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[32][12] ), .B2(n3832), .ZN(n3817) );
  INV_X1 U4845 ( .A(n3817), .ZN(\xmem_inst/n3478 ) );
  OAI22_X1 U4846 ( .A1(n3835), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[32][13] ), .B2(n3832), .ZN(n3818) );
  INV_X1 U4847 ( .A(n3818), .ZN(\xmem_inst/n3479 ) );
  OAI22_X1 U4848 ( .A1(n3835), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[32][14] ), .B2(n3832), .ZN(n3819) );
  INV_X1 U4849 ( .A(n3819), .ZN(\xmem_inst/n3480 ) );
  OAI22_X1 U4850 ( .A1(n3835), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[32][15] ), .B2(n3834), .ZN(n5168) );
  OAI22_X1 U4851 ( .A1(n3835), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[32][16] ), .B2(n3832), .ZN(n3820) );
  INV_X1 U4852 ( .A(n3820), .ZN(\xmem_inst/n3482 ) );
  OAI22_X1 U4853 ( .A1(n3835), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[32][17] ), .B2(n3832), .ZN(n3821) );
  INV_X1 U4854 ( .A(n3821), .ZN(\xmem_inst/n3483 ) );
  OAI22_X1 U4855 ( .A1(n3835), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[32][18] ), .B2(n3832), .ZN(n3822) );
  INV_X1 U4856 ( .A(n3822), .ZN(\xmem_inst/n3484 ) );
  OAI22_X1 U4857 ( .A1(n3835), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[32][19] ), .B2(n3834), .ZN(n5169) );
  OAI22_X1 U4858 ( .A1(n3835), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[32][20] ), .B2(n3832), .ZN(n3823) );
  INV_X1 U4859 ( .A(n3823), .ZN(\xmem_inst/n3486 ) );
  OAI22_X1 U4860 ( .A1(n3835), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[32][21] ), .B2(n3832), .ZN(n3824) );
  INV_X1 U4861 ( .A(n3824), .ZN(\xmem_inst/n3487 ) );
  OAI22_X1 U4862 ( .A1(n3835), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[32][22] ), .B2(n3834), .ZN(n3825) );
  INV_X1 U4863 ( .A(n3825), .ZN(\xmem_inst/n3488 ) );
  OAI22_X1 U4864 ( .A1(n3835), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[32][23] ), .B2(n3834), .ZN(n3826) );
  INV_X1 U4865 ( .A(n3826), .ZN(\xmem_inst/n3489 ) );
  OAI22_X1 U4866 ( .A1(n3835), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[32][24] ), .B2(n3834), .ZN(n3827) );
  INV_X1 U4867 ( .A(n3827), .ZN(\xmem_inst/n3490 ) );
  OAI22_X1 U4868 ( .A1(n3835), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[32][25] ), .B2(n3832), .ZN(n3828) );
  INV_X1 U4869 ( .A(n3828), .ZN(\xmem_inst/n3491 ) );
  OAI22_X1 U4870 ( .A1(n3835), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[32][26] ), .B2(n3834), .ZN(n3829) );
  INV_X1 U4871 ( .A(n3829), .ZN(\xmem_inst/n3492 ) );
  OAI22_X1 U4872 ( .A1(n3835), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[32][27] ), .B2(n3832), .ZN(n3830) );
  INV_X1 U4873 ( .A(n3830), .ZN(\xmem_inst/n3493 ) );
  OAI22_X1 U4874 ( .A1(n3835), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[32][28] ), .B2(n3834), .ZN(n3831) );
  INV_X1 U4875 ( .A(n3831), .ZN(\xmem_inst/n3494 ) );
  OAI22_X1 U4876 ( .A1(n3835), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[32][29] ), .B2(n3832), .ZN(n3833) );
  INV_X1 U4877 ( .A(n3833), .ZN(\xmem_inst/n3495 ) );
  OAI22_X1 U4878 ( .A1(n3835), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[32][30] ), .B2(n3834), .ZN(n5170) );
  OAI22_X1 U4879 ( .A1(n3835), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[32][31] ), .B2(n3834), .ZN(n5171) );
  NOR2_X2 U4880 ( .A1(n3933), .A2(n3890), .ZN(n3856) );
  INV_X2 U4881 ( .A(n3858), .ZN(n3859) );
  OAI22_X1 U4882 ( .A1(n3859), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[33][0] ), .B2(n3858), .ZN(n3836) );
  INV_X1 U4883 ( .A(n3836), .ZN(\xmem_inst/n3498 ) );
  OAI22_X1 U4884 ( .A1(n3859), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[33][1] ), .B2(n3856), .ZN(n3837) );
  INV_X1 U4885 ( .A(n3837), .ZN(\xmem_inst/n3499 ) );
  OAI22_X1 U4886 ( .A1(n3859), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[33][2] ), .B2(n3856), .ZN(n3838) );
  INV_X1 U4887 ( .A(n3838), .ZN(\xmem_inst/n3500 ) );
  OAI22_X1 U4888 ( .A1(n3859), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[33][3] ), .B2(n3856), .ZN(n3839) );
  INV_X1 U4889 ( .A(n3839), .ZN(\xmem_inst/n3501 ) );
  OAI22_X1 U4890 ( .A1(n3859), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[33][4] ), .B2(n3856), .ZN(n3840) );
  INV_X1 U4891 ( .A(n3840), .ZN(\xmem_inst/n3502 ) );
  OAI22_X1 U4892 ( .A1(n3859), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[33][5] ), .B2(n3856), .ZN(n3841) );
  INV_X1 U4893 ( .A(n3841), .ZN(\xmem_inst/n3503 ) );
  OAI22_X1 U4894 ( .A1(n3859), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[33][6] ), .B2(n3856), .ZN(n3842) );
  INV_X1 U4895 ( .A(n3842), .ZN(\xmem_inst/n3504 ) );
  OAI22_X1 U4896 ( .A1(n3859), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[33][7] ), .B2(n3856), .ZN(n3843) );
  INV_X1 U4897 ( .A(n3843), .ZN(\xmem_inst/n3505 ) );
  OAI22_X1 U4898 ( .A1(n3859), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[33][8] ), .B2(n3856), .ZN(n3844) );
  INV_X1 U4899 ( .A(n3844), .ZN(\xmem_inst/n3506 ) );
  OAI22_X1 U4900 ( .A1(n3859), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[33][9] ), .B2(n3856), .ZN(n3845) );
  INV_X1 U4901 ( .A(n3845), .ZN(\xmem_inst/n3507 ) );
  OAI22_X1 U4902 ( .A1(n3859), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[33][10] ), .B2(n3856), .ZN(n3846) );
  INV_X1 U4903 ( .A(n3846), .ZN(\xmem_inst/n3508 ) );
  OAI22_X1 U4904 ( .A1(n3859), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[33][11] ), .B2(n3856), .ZN(n3847) );
  INV_X1 U4905 ( .A(n3847), .ZN(\xmem_inst/n3509 ) );
  OAI22_X1 U4906 ( .A1(n3859), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[33][12] ), .B2(n3856), .ZN(n3848) );
  INV_X1 U4907 ( .A(n3848), .ZN(\xmem_inst/n3510 ) );
  OAI22_X1 U4908 ( .A1(n3859), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[33][13] ), .B2(n3856), .ZN(n3849) );
  INV_X1 U4909 ( .A(n3849), .ZN(\xmem_inst/n3511 ) );
  OAI22_X1 U4910 ( .A1(n3859), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[33][14] ), .B2(n3856), .ZN(n3850) );
  INV_X1 U4911 ( .A(n3850), .ZN(\xmem_inst/n3512 ) );
  OAI22_X1 U4912 ( .A1(n3859), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[33][15] ), .B2(n3858), .ZN(n5172) );
  OAI22_X1 U4913 ( .A1(n3859), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[33][16] ), .B2(n3856), .ZN(n3851) );
  INV_X1 U4914 ( .A(n3851), .ZN(\xmem_inst/n3514 ) );
  OAI22_X1 U4915 ( .A1(n3859), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[33][17] ), .B2(n3856), .ZN(n3852) );
  INV_X1 U4916 ( .A(n3852), .ZN(\xmem_inst/n3515 ) );
  OAI22_X1 U4917 ( .A1(n3859), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[33][18] ), .B2(n3856), .ZN(n3853) );
  INV_X1 U4918 ( .A(n3853), .ZN(\xmem_inst/n3516 ) );
  OAI22_X1 U4919 ( .A1(n3859), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[33][19] ), .B2(n3858), .ZN(n5173) );
  OAI22_X1 U4920 ( .A1(n3859), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[33][20] ), .B2(n3856), .ZN(n5174) );
  OAI22_X1 U4921 ( .A1(n3859), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[33][21] ), .B2(n3856), .ZN(n5175) );
  OAI22_X1 U4922 ( .A1(n3859), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[33][22] ), .B2(n3858), .ZN(n5176) );
  OAI22_X1 U4923 ( .A1(n3859), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[33][23] ), .B2(n3858), .ZN(n5177) );
  OAI22_X1 U4924 ( .A1(n3859), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[33][24] ), .B2(n3858), .ZN(n5178) );
  OAI22_X1 U4925 ( .A1(n3859), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[33][25] ), .B2(n3856), .ZN(n3854) );
  INV_X1 U4926 ( .A(n3854), .ZN(\xmem_inst/n3523 ) );
  OAI22_X1 U4927 ( .A1(n3859), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[33][26] ), .B2(n3858), .ZN(n5179) );
  OAI22_X1 U4928 ( .A1(n3859), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[33][27] ), .B2(n3856), .ZN(n3855) );
  INV_X1 U4929 ( .A(n3855), .ZN(\xmem_inst/n3525 ) );
  OAI22_X1 U4930 ( .A1(n3859), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[33][28] ), .B2(n3858), .ZN(n5180) );
  OAI22_X1 U4931 ( .A1(n3859), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[33][29] ), .B2(n3856), .ZN(n3857) );
  INV_X1 U4932 ( .A(n3857), .ZN(\xmem_inst/n3527 ) );
  OAI22_X1 U4933 ( .A1(n3859), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[33][30] ), .B2(n3858), .ZN(n5181) );
  OAI22_X1 U4934 ( .A1(n3859), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[33][31] ), .B2(n3858), .ZN(n5182) );
  NOR2_X2 U4935 ( .A1(n3970), .A2(n3890), .ZN(n3869) );
  INV_X2 U4936 ( .A(n3871), .ZN(n3872) );
  OAI22_X1 U4937 ( .A1(n3872), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[34][0] ), .B2(n3871), .ZN(n5183) );
  OAI22_X1 U4938 ( .A1(n3872), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[34][1] ), .B2(n3869), .ZN(n5184) );
  OAI22_X1 U4939 ( .A1(n3872), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[34][2] ), .B2(n3869), .ZN(n5185) );
  OAI22_X1 U4940 ( .A1(n3872), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[34][3] ), .B2(n3869), .ZN(n5186) );
  OAI22_X1 U4941 ( .A1(n3872), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[34][4] ), .B2(n3869), .ZN(n5187) );
  OAI22_X1 U4942 ( .A1(n3872), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[34][5] ), .B2(n3869), .ZN(n3860) );
  INV_X1 U4943 ( .A(n3860), .ZN(\xmem_inst/n3535 ) );
  OAI22_X1 U4944 ( .A1(n3872), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[34][6] ), .B2(n3869), .ZN(n3861) );
  INV_X1 U4945 ( .A(n3861), .ZN(\xmem_inst/n3536 ) );
  OAI22_X1 U4946 ( .A1(n3872), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[34][7] ), .B2(n3869), .ZN(n3862) );
  INV_X1 U4947 ( .A(n3862), .ZN(\xmem_inst/n3537 ) );
  OAI22_X1 U4948 ( .A1(n3872), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[34][8] ), .B2(n3869), .ZN(n3863) );
  INV_X1 U4949 ( .A(n3863), .ZN(\xmem_inst/n3538 ) );
  OAI22_X1 U4950 ( .A1(n3872), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[34][9] ), .B2(n3869), .ZN(n3864) );
  INV_X1 U4951 ( .A(n3864), .ZN(\xmem_inst/n3539 ) );
  OAI22_X1 U4952 ( .A1(n3872), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[34][10] ), .B2(n3869), .ZN(n5188) );
  OAI22_X1 U4953 ( .A1(n3872), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[34][11] ), .B2(n3869), .ZN(n3865) );
  INV_X1 U4954 ( .A(n3865), .ZN(\xmem_inst/n3541 ) );
  OAI22_X1 U4955 ( .A1(n3872), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[34][12] ), .B2(n3869), .ZN(n5189) );
  OAI22_X1 U4956 ( .A1(n3872), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[34][13] ), .B2(n3869), .ZN(n5190) );
  OAI22_X1 U4957 ( .A1(n3872), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[34][14] ), .B2(n3869), .ZN(n3866) );
  INV_X1 U4958 ( .A(n3866), .ZN(\xmem_inst/n3544 ) );
  OAI22_X1 U4959 ( .A1(n3872), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[34][15] ), .B2(n3871), .ZN(n5191) );
  OAI22_X1 U4960 ( .A1(n3872), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[34][16] ), .B2(n3869), .ZN(n5192) );
  OAI22_X1 U4961 ( .A1(n3872), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[34][17] ), .B2(n3869), .ZN(n5193) );
  OAI22_X1 U4962 ( .A1(n3872), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[34][18] ), .B2(n3869), .ZN(n5194) );
  OAI22_X1 U4963 ( .A1(n3872), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[34][19] ), .B2(n3871), .ZN(n5195) );
  OAI22_X1 U4964 ( .A1(n3872), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[34][20] ), .B2(n3869), .ZN(n5196) );
  OAI22_X1 U4965 ( .A1(n3872), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[34][21] ), .B2(n3869), .ZN(n5197) );
  OAI22_X1 U4966 ( .A1(n3872), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[34][22] ), .B2(n3871), .ZN(n5198) );
  OAI22_X1 U4967 ( .A1(n3872), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[34][23] ), .B2(n3871), .ZN(n5199) );
  OAI22_X1 U4968 ( .A1(n3872), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[34][24] ), .B2(n3871), .ZN(n5200) );
  OAI22_X1 U4969 ( .A1(n3872), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[34][25] ), .B2(n3869), .ZN(n3867) );
  INV_X1 U4970 ( .A(n3867), .ZN(\xmem_inst/n3555 ) );
  OAI22_X1 U4971 ( .A1(n3872), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[34][26] ), .B2(n3871), .ZN(n5201) );
  OAI22_X1 U4972 ( .A1(n3872), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[34][27] ), .B2(n3869), .ZN(n3868) );
  INV_X1 U4973 ( .A(n3868), .ZN(\xmem_inst/n3557 ) );
  OAI22_X1 U4974 ( .A1(n3872), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[34][28] ), .B2(n3871), .ZN(n5202) );
  OAI22_X1 U4975 ( .A1(n3872), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[34][29] ), .B2(n3869), .ZN(n3870) );
  INV_X1 U4976 ( .A(n3870), .ZN(\xmem_inst/n3559 ) );
  OAI22_X1 U4977 ( .A1(n3872), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[34][30] ), .B2(n3871), .ZN(n5203) );
  OAI22_X1 U4978 ( .A1(n3872), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[34][31] ), .B2(n3871), .ZN(n5204) );
  NOR2_X2 U4979 ( .A1(n3890), .A2(n3873), .ZN(n3876) );
  OAI22_X1 U4980 ( .A1(n3875), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[35][0] ), .B2(n3876), .ZN(n5205) );
  INV_X2 U4981 ( .A(n3877), .ZN(n3875) );
  OAI22_X1 U4982 ( .A1(n3875), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[35][1] ), .B2(n3876), .ZN(n5206) );
  OAI22_X1 U4983 ( .A1(n3875), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[35][2] ), .B2(n3876), .ZN(n5207) );
  OAI22_X1 U4984 ( .A1(n3875), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[35][3] ), .B2(n3876), .ZN(n5208) );
  OAI22_X1 U4985 ( .A1(n3875), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[35][4] ), .B2(n3876), .ZN(n5209) );
  OAI22_X1 U4986 ( .A1(n3875), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[35][5] ), .B2(n3876), .ZN(n5210) );
  OAI22_X1 U4987 ( .A1(n3875), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[35][6] ), .B2(n3876), .ZN(n5211) );
  OAI22_X1 U4988 ( .A1(n3875), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[35][7] ), .B2(n3876), .ZN(n5212) );
  OAI22_X1 U4989 ( .A1(n3875), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[35][8] ), .B2(n3876), .ZN(n5213) );
  OAI22_X1 U4990 ( .A1(n3875), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[35][9] ), .B2(n3876), .ZN(n5214) );
  OAI22_X1 U4991 ( .A1(n3875), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[35][10] ), .B2(n3876), .ZN(n5215) );
  OAI22_X1 U4992 ( .A1(n3875), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[35][11] ), .B2(n3876), .ZN(n5216) );
  OAI22_X1 U4993 ( .A1(n3875), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[35][12] ), .B2(n3877), .ZN(n3874) );
  INV_X1 U4994 ( .A(n3874), .ZN(\xmem_inst/n3574 ) );
  OAI22_X1 U4995 ( .A1(n3875), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[35][13] ), .B2(n3876), .ZN(n5217) );
  OAI22_X1 U4996 ( .A1(n3875), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[35][14] ), .B2(n3876), .ZN(n5218) );
  OAI22_X1 U4997 ( .A1(n3875), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[35][15] ), .B2(n3876), .ZN(n5219) );
  OAI22_X1 U4998 ( .A1(n3875), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[35][16] ), .B2(n3877), .ZN(n5220) );
  OAI22_X1 U4999 ( .A1(n3875), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[35][17] ), .B2(n3876), .ZN(n5221) );
  OAI22_X1 U5000 ( .A1(n3875), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[35][18] ), .B2(n3876), .ZN(n5222) );
  OAI22_X1 U5001 ( .A1(n3875), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[35][19] ), .B2(n3877), .ZN(n5223) );
  OAI22_X1 U5002 ( .A1(n3875), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[35][20] ), .B2(n3876), .ZN(n5224) );
  OAI22_X1 U5003 ( .A1(n3875), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[35][21] ), .B2(n3876), .ZN(n5225) );
  OAI22_X1 U5004 ( .A1(n3875), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[35][22] ), .B2(n3877), .ZN(n5226) );
  OAI22_X1 U5005 ( .A1(n3875), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[35][23] ), .B2(n3877), .ZN(n5227) );
  OAI22_X1 U5006 ( .A1(n3875), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[35][24] ), .B2(n3877), .ZN(n5228) );
  OAI22_X1 U5007 ( .A1(n3875), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[35][25] ), .B2(n3876), .ZN(n5229) );
  OAI22_X1 U5008 ( .A1(n3875), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[35][26] ), .B2(n3877), .ZN(n5230) );
  OAI22_X1 U5009 ( .A1(n3875), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[35][27] ), .B2(n3876), .ZN(n5231) );
  OAI22_X1 U5010 ( .A1(n3875), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[35][28] ), .B2(n3877), .ZN(n5232) );
  OAI22_X1 U5011 ( .A1(n3875), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[35][29] ), .B2(n3876), .ZN(n5233) );
  OAI22_X1 U5012 ( .A1(n3875), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[35][30] ), .B2(n3877), .ZN(n5234) );
  OAI22_X1 U5013 ( .A1(n3875), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[35][31] ), .B2(n3877), .ZN(n5235) );
  NOR2_X2 U5014 ( .A1(n3890), .A2(n3878), .ZN(n3879) );
  INV_X2 U5015 ( .A(n3880), .ZN(n3881) );
  OAI22_X1 U5016 ( .A1(n3881), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[36][0] ), .B2(n3880), .ZN(n5236) );
  OAI22_X1 U5017 ( .A1(n3881), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[36][1] ), .B2(n3879), .ZN(n5237) );
  OAI22_X1 U5018 ( .A1(n3881), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[36][2] ), .B2(n3879), .ZN(n5238) );
  OAI22_X1 U5019 ( .A1(n3881), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[36][3] ), .B2(n3879), .ZN(n5239) );
  OAI22_X1 U5020 ( .A1(n3881), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[36][4] ), .B2(n3879), .ZN(n5240) );
  OAI22_X1 U5021 ( .A1(n3881), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[36][5] ), .B2(n3879), .ZN(n5241) );
  OAI22_X1 U5022 ( .A1(n3881), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[36][6] ), .B2(n3879), .ZN(n5242) );
  OAI22_X1 U5023 ( .A1(n3881), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[36][7] ), .B2(n3879), .ZN(n5243) );
  OAI22_X1 U5024 ( .A1(n3881), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[36][8] ), .B2(n3879), .ZN(n5244) );
  OAI22_X1 U5025 ( .A1(n3881), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[36][9] ), .B2(n3879), .ZN(n5245) );
  OAI22_X1 U5026 ( .A1(n3881), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[36][10] ), .B2(n3879), .ZN(n5246) );
  OAI22_X1 U5027 ( .A1(n3881), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[36][11] ), .B2(n3879), .ZN(n5247) );
  OAI22_X1 U5028 ( .A1(n3881), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[36][12] ), .B2(n3879), .ZN(n5248) );
  OAI22_X1 U5029 ( .A1(n3881), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[36][13] ), .B2(n3879), .ZN(n5249) );
  OAI22_X1 U5030 ( .A1(n3881), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[36][14] ), .B2(n3879), .ZN(n5250) );
  OAI22_X1 U5031 ( .A1(n3881), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[36][15] ), .B2(n3879), .ZN(n5251) );
  OAI22_X1 U5032 ( .A1(n3881), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[36][16] ), .B2(n3880), .ZN(n5252) );
  OAI22_X1 U5033 ( .A1(n3881), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[36][17] ), .B2(n3879), .ZN(n5253) );
  OAI22_X1 U5034 ( .A1(n3881), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[36][18] ), .B2(n3879), .ZN(n5254) );
  OAI22_X1 U5035 ( .A1(n3881), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[36][19] ), .B2(n3880), .ZN(n5255) );
  OAI22_X1 U5036 ( .A1(n3881), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[36][20] ), .B2(n3879), .ZN(n5256) );
  OAI22_X1 U5037 ( .A1(n3881), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[36][21] ), .B2(n3879), .ZN(n5257) );
  OAI22_X1 U5038 ( .A1(n3881), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[36][22] ), .B2(n3880), .ZN(n5258) );
  OAI22_X1 U5039 ( .A1(n3881), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[36][23] ), .B2(n3880), .ZN(n5259) );
  OAI22_X1 U5040 ( .A1(n3881), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[36][24] ), .B2(n3880), .ZN(n5260) );
  OAI22_X1 U5041 ( .A1(n3881), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[36][25] ), .B2(n3879), .ZN(n5261) );
  OAI22_X1 U5042 ( .A1(n3881), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[36][26] ), .B2(n3880), .ZN(n5262) );
  OAI22_X1 U5043 ( .A1(n3881), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[36][27] ), .B2(n3879), .ZN(n5263) );
  OAI22_X1 U5044 ( .A1(n3881), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[36][28] ), .B2(n3880), .ZN(n5264) );
  OAI22_X1 U5045 ( .A1(n3881), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[36][29] ), .B2(n3879), .ZN(n5265) );
  OAI22_X1 U5046 ( .A1(n3881), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[36][30] ), .B2(n3880), .ZN(n5266) );
  OAI22_X1 U5047 ( .A1(n3881), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[36][31] ), .B2(n3880), .ZN(n5267) );
  NOR2_X2 U5048 ( .A1(n3890), .A2(n3882), .ZN(n3883) );
  INV_X2 U5049 ( .A(n3884), .ZN(n3885) );
  OAI22_X1 U5050 ( .A1(n3885), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[37][0] ), .B2(n3884), .ZN(n5268) );
  OAI22_X1 U5051 ( .A1(n3885), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[37][1] ), .B2(n3883), .ZN(n5269) );
  OAI22_X1 U5052 ( .A1(n3885), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[37][2] ), .B2(n3883), .ZN(n5270) );
  OAI22_X1 U5053 ( .A1(n3885), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[37][3] ), .B2(n3883), .ZN(n5271) );
  OAI22_X1 U5054 ( .A1(n3885), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[37][4] ), .B2(n3883), .ZN(n5272) );
  OAI22_X1 U5055 ( .A1(n3885), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[37][5] ), .B2(n3883), .ZN(n5273) );
  OAI22_X1 U5056 ( .A1(n3885), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[37][6] ), .B2(n3883), .ZN(n5274) );
  OAI22_X1 U5057 ( .A1(n3885), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[37][7] ), .B2(n3883), .ZN(n5275) );
  OAI22_X1 U5058 ( .A1(n3885), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[37][8] ), .B2(n3883), .ZN(n5276) );
  OAI22_X1 U5059 ( .A1(n3885), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[37][9] ), .B2(n3883), .ZN(n5277) );
  OAI22_X1 U5060 ( .A1(n3885), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[37][10] ), .B2(n3883), .ZN(n5278) );
  OAI22_X1 U5061 ( .A1(n3885), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[37][11] ), .B2(n3883), .ZN(n5279) );
  OAI22_X1 U5062 ( .A1(n3885), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[37][12] ), .B2(n3883), .ZN(n5280) );
  OAI22_X1 U5063 ( .A1(n3885), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[37][13] ), .B2(n3883), .ZN(n5281) );
  OAI22_X1 U5064 ( .A1(n3885), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[37][14] ), .B2(n3883), .ZN(n5282) );
  OAI22_X1 U5065 ( .A1(n3885), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[37][15] ), .B2(n3883), .ZN(n5283) );
  OAI22_X1 U5066 ( .A1(n3885), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[37][16] ), .B2(n3884), .ZN(n5284) );
  OAI22_X1 U5067 ( .A1(n3885), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[37][17] ), .B2(n3883), .ZN(n5285) );
  OAI22_X1 U5068 ( .A1(n3885), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[37][18] ), .B2(n3883), .ZN(n5286) );
  OAI22_X1 U5069 ( .A1(n3885), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[37][19] ), .B2(n3884), .ZN(n5287) );
  OAI22_X1 U5070 ( .A1(n3885), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[37][20] ), .B2(n3883), .ZN(n5288) );
  OAI22_X1 U5071 ( .A1(n3885), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[37][21] ), .B2(n3883), .ZN(n5289) );
  OAI22_X1 U5072 ( .A1(n3885), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[37][22] ), .B2(n3884), .ZN(n5290) );
  OAI22_X1 U5073 ( .A1(n3885), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[37][23] ), .B2(n3884), .ZN(n5291) );
  OAI22_X1 U5074 ( .A1(n3885), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[37][24] ), .B2(n3884), .ZN(n5292) );
  OAI22_X1 U5075 ( .A1(n3885), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[37][25] ), .B2(n3883), .ZN(n5293) );
  OAI22_X1 U5076 ( .A1(n3885), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[37][26] ), .B2(n3884), .ZN(n5294) );
  OAI22_X1 U5077 ( .A1(n3885), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[37][27] ), .B2(n3883), .ZN(n5295) );
  OAI22_X1 U5078 ( .A1(n3885), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[37][28] ), .B2(n3884), .ZN(n5296) );
  OAI22_X1 U5079 ( .A1(n3885), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[37][29] ), .B2(n3883), .ZN(n5297) );
  OAI22_X1 U5080 ( .A1(n3885), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[37][30] ), .B2(n3884), .ZN(n5298) );
  OAI22_X1 U5081 ( .A1(n3885), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[37][31] ), .B2(n3884), .ZN(n5299) );
  NOR2_X2 U5082 ( .A1(n3890), .A2(n3886), .ZN(n3887) );
  INV_X2 U5083 ( .A(n3888), .ZN(n3889) );
  OAI22_X1 U5084 ( .A1(n3889), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[38][0] ), .B2(n3888), .ZN(n5300) );
  OAI22_X1 U5085 ( .A1(n3889), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[38][1] ), .B2(n3887), .ZN(n5301) );
  OAI22_X1 U5086 ( .A1(n3889), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[38][2] ), .B2(n3887), .ZN(n5302) );
  OAI22_X1 U5087 ( .A1(n3889), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[38][3] ), .B2(n3887), .ZN(n5303) );
  OAI22_X1 U5088 ( .A1(n3889), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[38][4] ), .B2(n3887), .ZN(n5304) );
  OAI22_X1 U5089 ( .A1(n3889), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[38][5] ), .B2(n3887), .ZN(n5305) );
  OAI22_X1 U5090 ( .A1(n3889), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[38][6] ), .B2(n3887), .ZN(n5306) );
  OAI22_X1 U5091 ( .A1(n3889), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[38][7] ), .B2(n3887), .ZN(n5307) );
  OAI22_X1 U5092 ( .A1(n3889), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[38][8] ), .B2(n3887), .ZN(n5308) );
  OAI22_X1 U5093 ( .A1(n3889), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[38][9] ), .B2(n3887), .ZN(n5309) );
  OAI22_X1 U5094 ( .A1(n3889), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[38][10] ), .B2(n3887), .ZN(n5310) );
  OAI22_X1 U5095 ( .A1(n3889), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[38][11] ), .B2(n3887), .ZN(n5311) );
  OAI22_X1 U5096 ( .A1(n3889), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[38][12] ), .B2(n3887), .ZN(n5312) );
  OAI22_X1 U5097 ( .A1(n3889), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[38][13] ), .B2(n3887), .ZN(n5313) );
  OAI22_X1 U5098 ( .A1(n3889), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[38][14] ), .B2(n3887), .ZN(n5314) );
  OAI22_X1 U5099 ( .A1(n3889), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[38][15] ), .B2(n3887), .ZN(n5315) );
  OAI22_X1 U5100 ( .A1(n3889), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[38][16] ), .B2(n3888), .ZN(n5316) );
  OAI22_X1 U5101 ( .A1(n3889), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[38][17] ), .B2(n3887), .ZN(n5317) );
  OAI22_X1 U5102 ( .A1(n3889), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[38][18] ), .B2(n3887), .ZN(n5318) );
  OAI22_X1 U5103 ( .A1(n3889), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[38][19] ), .B2(n3888), .ZN(n5319) );
  OAI22_X1 U5104 ( .A1(n3889), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[38][20] ), .B2(n3887), .ZN(n5320) );
  OAI22_X1 U5105 ( .A1(n3889), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[38][21] ), .B2(n3887), .ZN(n5321) );
  OAI22_X1 U5106 ( .A1(n3889), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[38][22] ), .B2(n3888), .ZN(n5322) );
  OAI22_X1 U5107 ( .A1(n3889), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[38][23] ), .B2(n3888), .ZN(n5323) );
  OAI22_X1 U5108 ( .A1(n3889), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[38][24] ), .B2(n3888), .ZN(n5324) );
  OAI22_X1 U5109 ( .A1(n3889), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[38][25] ), .B2(n3887), .ZN(n5325) );
  OAI22_X1 U5110 ( .A1(n3889), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[38][26] ), .B2(n3888), .ZN(n5326) );
  OAI22_X1 U5111 ( .A1(n3889), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[38][27] ), .B2(n3887), .ZN(n5327) );
  OAI22_X1 U5112 ( .A1(n3889), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[38][28] ), .B2(n3888), .ZN(n5328) );
  OAI22_X1 U5113 ( .A1(n3889), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[38][29] ), .B2(n3887), .ZN(n5329) );
  OAI22_X1 U5114 ( .A1(n3889), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[38][30] ), .B2(n3888), .ZN(n5330) );
  OAI22_X1 U5115 ( .A1(n3889), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[38][31] ), .B2(n3888), .ZN(n5331) );
  NOR2_X2 U5116 ( .A1(n3891), .A2(n3890), .ZN(n3893) );
  INV_X2 U5117 ( .A(n3894), .ZN(n3895) );
  OAI22_X1 U5118 ( .A1(n3895), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[39][0] ), .B2(n3893), .ZN(n5332) );
  OAI22_X1 U5119 ( .A1(n3895), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[39][1] ), .B2(n3893), .ZN(n5333) );
  OAI22_X1 U5120 ( .A1(n3895), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[39][2] ), .B2(n3893), .ZN(n5334) );
  OAI22_X1 U5121 ( .A1(n3895), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[39][3] ), .B2(n3893), .ZN(n5335) );
  OAI22_X1 U5122 ( .A1(n3895), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[39][4] ), .B2(n3894), .ZN(n3892) );
  INV_X1 U5123 ( .A(n3892), .ZN(\xmem_inst/n3694 ) );
  OAI22_X1 U5124 ( .A1(n3895), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[39][5] ), .B2(n3893), .ZN(n5336) );
  OAI22_X1 U5125 ( .A1(n3895), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[39][6] ), .B2(n3893), .ZN(n5337) );
  OAI22_X1 U5126 ( .A1(n3895), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[39][7] ), .B2(n3893), .ZN(n5338) );
  OAI22_X1 U5127 ( .A1(n3895), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[39][8] ), .B2(n3893), .ZN(n5339) );
  OAI22_X1 U5128 ( .A1(n3895), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[39][9] ), .B2(n3893), .ZN(n5340) );
  OAI22_X1 U5129 ( .A1(n3895), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[39][10] ), .B2(n3893), .ZN(n5341) );
  OAI22_X1 U5130 ( .A1(n3895), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[39][11] ), .B2(n3893), .ZN(n5342) );
  OAI22_X1 U5131 ( .A1(n3895), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[39][12] ), .B2(n3893), .ZN(n5343) );
  OAI22_X1 U5132 ( .A1(n3895), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[39][13] ), .B2(n3893), .ZN(n5344) );
  OAI22_X1 U5133 ( .A1(n3895), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[39][14] ), .B2(n3893), .ZN(n5345) );
  OAI22_X1 U5134 ( .A1(n3895), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[39][15] ), .B2(n3894), .ZN(n5346) );
  OAI22_X1 U5135 ( .A1(n3895), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[39][16] ), .B2(n3893), .ZN(n5347) );
  OAI22_X1 U5136 ( .A1(n3895), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[39][17] ), .B2(n3893), .ZN(n5348) );
  OAI22_X1 U5137 ( .A1(n3895), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[39][18] ), .B2(n3893), .ZN(n5349) );
  OAI22_X1 U5138 ( .A1(n3895), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[39][19] ), .B2(n3894), .ZN(n5350) );
  OAI22_X1 U5139 ( .A1(n3895), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[39][20] ), .B2(n3893), .ZN(n5351) );
  OAI22_X1 U5140 ( .A1(n3895), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[39][21] ), .B2(n3893), .ZN(n5352) );
  OAI22_X1 U5141 ( .A1(n3895), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[39][22] ), .B2(n3894), .ZN(n5353) );
  OAI22_X1 U5142 ( .A1(n3895), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[39][23] ), .B2(n3894), .ZN(n5354) );
  OAI22_X1 U5143 ( .A1(n3895), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[39][24] ), .B2(n3894), .ZN(n5355) );
  OAI22_X1 U5144 ( .A1(n3895), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[39][25] ), .B2(n3893), .ZN(n5356) );
  OAI22_X1 U5145 ( .A1(n3895), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[39][26] ), .B2(n3894), .ZN(n5357) );
  OAI22_X1 U5146 ( .A1(n3895), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[39][27] ), .B2(n3893), .ZN(n5358) );
  OAI22_X1 U5147 ( .A1(n3895), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[39][28] ), .B2(n3894), .ZN(n5359) );
  OAI22_X1 U5148 ( .A1(n3895), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[39][29] ), .B2(n3893), .ZN(n5360) );
  OAI22_X1 U5149 ( .A1(n3895), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[39][30] ), .B2(n3894), .ZN(n5361) );
  OAI22_X1 U5150 ( .A1(n3895), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[39][31] ), .B2(n3894), .ZN(n5362) );
  NAND4_X1 U5151 ( .A1(xmem_addr[5]), .A2(xmem_addr[3]), .A3(n3896), .A4(n4081), .ZN(n3969) );
  NOR2_X2 U5152 ( .A1(n3969), .A2(n3897), .ZN(n3927) );
  INV_X2 U5153 ( .A(n3930), .ZN(n3931) );
  OAI22_X1 U5154 ( .A1(n3931), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[40][0] ), .B2(n3930), .ZN(n3898) );
  INV_X1 U5155 ( .A(n3898), .ZN(\xmem_inst/n3722 ) );
  OAI22_X1 U5156 ( .A1(n3931), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[40][1] ), .B2(n3927), .ZN(n3899) );
  INV_X1 U5157 ( .A(n3899), .ZN(\xmem_inst/n3723 ) );
  OAI22_X1 U5158 ( .A1(n3931), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[40][2] ), .B2(n3927), .ZN(n3900) );
  INV_X1 U5159 ( .A(n3900), .ZN(\xmem_inst/n3724 ) );
  OAI22_X1 U5160 ( .A1(n3931), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[40][3] ), .B2(n3927), .ZN(n3901) );
  INV_X1 U5161 ( .A(n3901), .ZN(\xmem_inst/n3725 ) );
  OAI22_X1 U5162 ( .A1(n3931), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[40][4] ), .B2(n3927), .ZN(n3902) );
  INV_X1 U5163 ( .A(n3902), .ZN(\xmem_inst/n3726 ) );
  OAI22_X1 U5164 ( .A1(n3931), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[40][5] ), .B2(n3927), .ZN(n3903) );
  INV_X1 U5165 ( .A(n3903), .ZN(\xmem_inst/n3727 ) );
  OAI22_X1 U5166 ( .A1(n3931), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[40][6] ), .B2(n3927), .ZN(n3904) );
  INV_X1 U5167 ( .A(n3904), .ZN(\xmem_inst/n3728 ) );
  OAI22_X1 U5168 ( .A1(n3931), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[40][7] ), .B2(n3927), .ZN(n3905) );
  INV_X1 U5169 ( .A(n3905), .ZN(\xmem_inst/n3729 ) );
  OAI22_X1 U5170 ( .A1(n3931), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[40][8] ), .B2(n3927), .ZN(n3906) );
  INV_X1 U5171 ( .A(n3906), .ZN(\xmem_inst/n3730 ) );
  OAI22_X1 U5172 ( .A1(n3931), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[40][9] ), .B2(n3927), .ZN(n3907) );
  INV_X1 U5173 ( .A(n3907), .ZN(\xmem_inst/n3731 ) );
  OAI22_X1 U5174 ( .A1(n3931), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[40][10] ), .B2(n3927), .ZN(n3908) );
  INV_X1 U5175 ( .A(n3908), .ZN(\xmem_inst/n3732 ) );
  OAI22_X1 U5176 ( .A1(n3931), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[40][11] ), .B2(n3927), .ZN(n3909) );
  INV_X1 U5177 ( .A(n3909), .ZN(\xmem_inst/n3733 ) );
  OAI22_X1 U5178 ( .A1(n3931), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[40][12] ), .B2(n3927), .ZN(n3910) );
  INV_X1 U5179 ( .A(n3910), .ZN(\xmem_inst/n3734 ) );
  OAI22_X1 U5180 ( .A1(n3931), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[40][13] ), .B2(n3927), .ZN(n3911) );
  INV_X1 U5181 ( .A(n3911), .ZN(\xmem_inst/n3735 ) );
  OAI22_X1 U5182 ( .A1(n3931), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[40][14] ), .B2(n3927), .ZN(n3912) );
  INV_X1 U5183 ( .A(n3912), .ZN(\xmem_inst/n3736 ) );
  OAI22_X1 U5184 ( .A1(n3931), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[40][15] ), .B2(n3930), .ZN(n3913) );
  INV_X1 U5185 ( .A(n3913), .ZN(\xmem_inst/n3737 ) );
  OAI22_X1 U5186 ( .A1(n3931), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[40][16] ), .B2(n3927), .ZN(n3914) );
  INV_X1 U5187 ( .A(n3914), .ZN(\xmem_inst/n3738 ) );
  OAI22_X1 U5188 ( .A1(n3931), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[40][17] ), .B2(n3927), .ZN(n3915) );
  INV_X1 U5189 ( .A(n3915), .ZN(\xmem_inst/n3739 ) );
  OAI22_X1 U5190 ( .A1(n3931), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[40][18] ), .B2(n3927), .ZN(n3916) );
  INV_X1 U5191 ( .A(n3916), .ZN(\xmem_inst/n3740 ) );
  OAI22_X1 U5192 ( .A1(n3931), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[40][19] ), .B2(n3930), .ZN(n3917) );
  INV_X1 U5193 ( .A(n3917), .ZN(\xmem_inst/n3741 ) );
  OAI22_X1 U5194 ( .A1(n3931), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[40][20] ), .B2(n3927), .ZN(n3918) );
  INV_X1 U5195 ( .A(n3918), .ZN(\xmem_inst/n3742 ) );
  OAI22_X1 U5196 ( .A1(n3931), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[40][21] ), .B2(n3927), .ZN(n3919) );
  INV_X1 U5197 ( .A(n3919), .ZN(\xmem_inst/n3743 ) );
  OAI22_X1 U5198 ( .A1(n3931), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[40][22] ), .B2(n3930), .ZN(n3920) );
  INV_X1 U5199 ( .A(n3920), .ZN(\xmem_inst/n3744 ) );
  OAI22_X1 U5200 ( .A1(n3931), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[40][23] ), .B2(n3930), .ZN(n3921) );
  INV_X1 U5201 ( .A(n3921), .ZN(\xmem_inst/n3745 ) );
  OAI22_X1 U5202 ( .A1(n3931), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[40][24] ), .B2(n3930), .ZN(n3922) );
  INV_X1 U5203 ( .A(n3922), .ZN(\xmem_inst/n3746 ) );
  OAI22_X1 U5204 ( .A1(n3931), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[40][25] ), .B2(n3927), .ZN(n3923) );
  INV_X1 U5205 ( .A(n3923), .ZN(\xmem_inst/n3747 ) );
  OAI22_X1 U5206 ( .A1(n3931), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[40][26] ), .B2(n3930), .ZN(n3924) );
  INV_X1 U5207 ( .A(n3924), .ZN(\xmem_inst/n3748 ) );
  OAI22_X1 U5208 ( .A1(n3931), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[40][27] ), .B2(n3927), .ZN(n3925) );
  INV_X1 U5209 ( .A(n3925), .ZN(\xmem_inst/n3749 ) );
  OAI22_X1 U5210 ( .A1(n3931), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[40][28] ), .B2(n3930), .ZN(n3926) );
  INV_X1 U5211 ( .A(n3926), .ZN(\xmem_inst/n3750 ) );
  OAI22_X1 U5212 ( .A1(n3931), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[40][29] ), .B2(n3927), .ZN(n3928) );
  INV_X1 U5213 ( .A(n3928), .ZN(\xmem_inst/n3751 ) );
  OAI22_X1 U5214 ( .A1(n3931), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[40][30] ), .B2(n3930), .ZN(n3929) );
  INV_X1 U5215 ( .A(n3929), .ZN(\xmem_inst/n3752 ) );
  OAI22_X1 U5216 ( .A1(n3931), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[40][31] ), .B2(n3930), .ZN(n3932) );
  INV_X1 U5217 ( .A(n3932), .ZN(\xmem_inst/n3753 ) );
  NOR2_X2 U5218 ( .A1(n3969), .A2(n3933), .ZN(n3963) );
  INV_X2 U5219 ( .A(n3966), .ZN(n3967) );
  OAI22_X1 U5220 ( .A1(n3967), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[41][0] ), .B2(n3966), .ZN(n3934) );
  INV_X1 U5221 ( .A(n3934), .ZN(\xmem_inst/n3754 ) );
  OAI22_X1 U5222 ( .A1(n3967), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[41][1] ), .B2(n3963), .ZN(n3935) );
  INV_X1 U5223 ( .A(n3935), .ZN(\xmem_inst/n3755 ) );
  OAI22_X1 U5224 ( .A1(n3967), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[41][2] ), .B2(n3963), .ZN(n3936) );
  INV_X1 U5225 ( .A(n3936), .ZN(\xmem_inst/n3756 ) );
  OAI22_X1 U5226 ( .A1(n3967), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[41][3] ), .B2(n3963), .ZN(n3937) );
  INV_X1 U5227 ( .A(n3937), .ZN(\xmem_inst/n3757 ) );
  OAI22_X1 U5228 ( .A1(n3967), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[41][4] ), .B2(n3963), .ZN(n3938) );
  INV_X1 U5229 ( .A(n3938), .ZN(\xmem_inst/n3758 ) );
  OAI22_X1 U5230 ( .A1(n3967), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[41][5] ), .B2(n3963), .ZN(n3939) );
  INV_X1 U5231 ( .A(n3939), .ZN(\xmem_inst/n3759 ) );
  OAI22_X1 U5232 ( .A1(n3967), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[41][6] ), .B2(n3963), .ZN(n3940) );
  INV_X1 U5233 ( .A(n3940), .ZN(\xmem_inst/n3760 ) );
  OAI22_X1 U5234 ( .A1(n3967), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[41][7] ), .B2(n3963), .ZN(n3941) );
  INV_X1 U5235 ( .A(n3941), .ZN(\xmem_inst/n3761 ) );
  OAI22_X1 U5236 ( .A1(n3967), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[41][8] ), .B2(n3963), .ZN(n3942) );
  INV_X1 U5237 ( .A(n3942), .ZN(\xmem_inst/n3762 ) );
  OAI22_X1 U5238 ( .A1(n3967), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[41][9] ), .B2(n3963), .ZN(n3943) );
  INV_X1 U5239 ( .A(n3943), .ZN(\xmem_inst/n3763 ) );
  OAI22_X1 U5240 ( .A1(n3967), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[41][10] ), .B2(n3963), .ZN(n3944) );
  INV_X1 U5241 ( .A(n3944), .ZN(\xmem_inst/n3764 ) );
  OAI22_X1 U5242 ( .A1(n3967), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[41][11] ), .B2(n3963), .ZN(n3945) );
  INV_X1 U5243 ( .A(n3945), .ZN(\xmem_inst/n3765 ) );
  OAI22_X1 U5244 ( .A1(n3967), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[41][12] ), .B2(n3963), .ZN(n3946) );
  INV_X1 U5245 ( .A(n3946), .ZN(\xmem_inst/n3766 ) );
  OAI22_X1 U5246 ( .A1(n3967), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[41][13] ), .B2(n3963), .ZN(n3947) );
  INV_X1 U5247 ( .A(n3947), .ZN(\xmem_inst/n3767 ) );
  OAI22_X1 U5248 ( .A1(n3967), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[41][14] ), .B2(n3963), .ZN(n3948) );
  INV_X1 U5249 ( .A(n3948), .ZN(\xmem_inst/n3768 ) );
  OAI22_X1 U5250 ( .A1(n3967), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[41][15] ), .B2(n3966), .ZN(n3949) );
  INV_X1 U5251 ( .A(n3949), .ZN(\xmem_inst/n3769 ) );
  OAI22_X1 U5252 ( .A1(n3967), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[41][16] ), .B2(n3963), .ZN(n3950) );
  INV_X1 U5253 ( .A(n3950), .ZN(\xmem_inst/n3770 ) );
  OAI22_X1 U5254 ( .A1(n3967), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[41][17] ), .B2(n3963), .ZN(n3951) );
  INV_X1 U5255 ( .A(n3951), .ZN(\xmem_inst/n3771 ) );
  OAI22_X1 U5256 ( .A1(n3967), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[41][18] ), .B2(n3963), .ZN(n3952) );
  INV_X1 U5257 ( .A(n3952), .ZN(\xmem_inst/n3772 ) );
  OAI22_X1 U5258 ( .A1(n3967), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[41][19] ), .B2(n3966), .ZN(n3953) );
  INV_X1 U5259 ( .A(n3953), .ZN(\xmem_inst/n3773 ) );
  OAI22_X1 U5260 ( .A1(n3967), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[41][20] ), .B2(n3963), .ZN(n3954) );
  INV_X1 U5261 ( .A(n3954), .ZN(\xmem_inst/n3774 ) );
  OAI22_X1 U5262 ( .A1(n3967), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[41][21] ), .B2(n3963), .ZN(n3955) );
  INV_X1 U5263 ( .A(n3955), .ZN(\xmem_inst/n3775 ) );
  OAI22_X1 U5264 ( .A1(n3967), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[41][22] ), .B2(n3966), .ZN(n3956) );
  INV_X1 U5265 ( .A(n3956), .ZN(\xmem_inst/n3776 ) );
  OAI22_X1 U5266 ( .A1(n3967), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[41][23] ), .B2(n3966), .ZN(n3957) );
  INV_X1 U5267 ( .A(n3957), .ZN(\xmem_inst/n3777 ) );
  OAI22_X1 U5268 ( .A1(n3967), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[41][24] ), .B2(n3966), .ZN(n3958) );
  INV_X1 U5269 ( .A(n3958), .ZN(\xmem_inst/n3778 ) );
  OAI22_X1 U5270 ( .A1(n3967), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[41][25] ), .B2(n3963), .ZN(n3959) );
  INV_X1 U5271 ( .A(n3959), .ZN(\xmem_inst/n3779 ) );
  OAI22_X1 U5272 ( .A1(n3967), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[41][26] ), .B2(n3966), .ZN(n3960) );
  INV_X1 U5273 ( .A(n3960), .ZN(\xmem_inst/n3780 ) );
  OAI22_X1 U5274 ( .A1(n3967), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[41][27] ), .B2(n3963), .ZN(n3961) );
  INV_X1 U5275 ( .A(n3961), .ZN(\xmem_inst/n3781 ) );
  OAI22_X1 U5276 ( .A1(n3967), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[41][28] ), .B2(n3966), .ZN(n3962) );
  INV_X1 U5277 ( .A(n3962), .ZN(\xmem_inst/n3782 ) );
  OAI22_X1 U5278 ( .A1(n3967), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[41][29] ), .B2(n3963), .ZN(n3964) );
  INV_X1 U5279 ( .A(n3964), .ZN(\xmem_inst/n3783 ) );
  OAI22_X1 U5280 ( .A1(n3967), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[41][30] ), .B2(n3966), .ZN(n3965) );
  INV_X1 U5281 ( .A(n3965), .ZN(\xmem_inst/n3784 ) );
  OAI22_X1 U5282 ( .A1(n3967), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[41][31] ), .B2(n3966), .ZN(n3968) );
  INV_X1 U5283 ( .A(n3968), .ZN(\xmem_inst/n3785 ) );
  NOR2_X2 U5284 ( .A1(n3970), .A2(n3969), .ZN(n4000) );
  INV_X2 U5285 ( .A(n4003), .ZN(n4004) );
  OAI22_X1 U5286 ( .A1(n4004), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[42][0] ), .B2(n4003), .ZN(n3971) );
  INV_X1 U5287 ( .A(n3971), .ZN(\xmem_inst/n3786 ) );
  OAI22_X1 U5288 ( .A1(n4004), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[42][1] ), .B2(n4000), .ZN(n3972) );
  INV_X1 U5289 ( .A(n3972), .ZN(\xmem_inst/n3787 ) );
  OAI22_X1 U5290 ( .A1(n4004), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[42][2] ), .B2(n4000), .ZN(n3973) );
  INV_X1 U5291 ( .A(n3973), .ZN(\xmem_inst/n3788 ) );
  OAI22_X1 U5292 ( .A1(n4004), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[42][3] ), .B2(n4000), .ZN(n3974) );
  INV_X1 U5293 ( .A(n3974), .ZN(\xmem_inst/n3789 ) );
  OAI22_X1 U5294 ( .A1(n4004), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[42][4] ), .B2(n4000), .ZN(n3975) );
  INV_X1 U5295 ( .A(n3975), .ZN(\xmem_inst/n3790 ) );
  OAI22_X1 U5296 ( .A1(n4004), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[42][5] ), .B2(n4000), .ZN(n3976) );
  INV_X1 U5297 ( .A(n3976), .ZN(\xmem_inst/n3791 ) );
  OAI22_X1 U5298 ( .A1(n4004), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[42][6] ), .B2(n4000), .ZN(n3977) );
  INV_X1 U5299 ( .A(n3977), .ZN(\xmem_inst/n3792 ) );
  OAI22_X1 U5300 ( .A1(n4004), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[42][7] ), .B2(n4000), .ZN(n3978) );
  INV_X1 U5301 ( .A(n3978), .ZN(\xmem_inst/n3793 ) );
  OAI22_X1 U5302 ( .A1(n4004), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[42][8] ), .B2(n4000), .ZN(n3979) );
  INV_X1 U5303 ( .A(n3979), .ZN(\xmem_inst/n3794 ) );
  OAI22_X1 U5304 ( .A1(n4004), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[42][9] ), .B2(n4000), .ZN(n3980) );
  INV_X1 U5305 ( .A(n3980), .ZN(\xmem_inst/n3795 ) );
  OAI22_X1 U5306 ( .A1(n4004), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[42][10] ), .B2(n4000), .ZN(n3981) );
  INV_X1 U5307 ( .A(n3981), .ZN(\xmem_inst/n3796 ) );
  OAI22_X1 U5308 ( .A1(n4004), .A2(s_data_in_x[11]), .B1(
        \xmem_inst/mem[42][11] ), .B2(n4000), .ZN(n3982) );
  INV_X1 U5309 ( .A(n3982), .ZN(\xmem_inst/n3797 ) );
  OAI22_X1 U5310 ( .A1(n4004), .A2(s_data_in_x[12]), .B1(
        \xmem_inst/mem[42][12] ), .B2(n4000), .ZN(n3983) );
  INV_X1 U5311 ( .A(n3983), .ZN(\xmem_inst/n3798 ) );
  OAI22_X1 U5312 ( .A1(n4004), .A2(s_data_in_x[13]), .B1(
        \xmem_inst/mem[42][13] ), .B2(n4000), .ZN(n3984) );
  INV_X1 U5313 ( .A(n3984), .ZN(\xmem_inst/n3799 ) );
  OAI22_X1 U5314 ( .A1(n4004), .A2(s_data_in_x[14]), .B1(
        \xmem_inst/mem[42][14] ), .B2(n4000), .ZN(n3985) );
  INV_X1 U5315 ( .A(n3985), .ZN(\xmem_inst/n3800 ) );
  OAI22_X1 U5316 ( .A1(n4004), .A2(s_data_in_x[15]), .B1(
        \xmem_inst/mem[42][15] ), .B2(n4003), .ZN(n3986) );
  INV_X1 U5317 ( .A(n3986), .ZN(\xmem_inst/n3801 ) );
  OAI22_X1 U5318 ( .A1(n4004), .A2(s_data_in_x[16]), .B1(
        \xmem_inst/mem[42][16] ), .B2(n4000), .ZN(n3987) );
  INV_X1 U5319 ( .A(n3987), .ZN(\xmem_inst/n3802 ) );
  OAI22_X1 U5320 ( .A1(n4004), .A2(s_data_in_x[17]), .B1(
        \xmem_inst/mem[42][17] ), .B2(n4000), .ZN(n3988) );
  INV_X1 U5321 ( .A(n3988), .ZN(\xmem_inst/n3803 ) );
  OAI22_X1 U5322 ( .A1(n4004), .A2(s_data_in_x[18]), .B1(
        \xmem_inst/mem[42][18] ), .B2(n4000), .ZN(n3989) );
  INV_X1 U5323 ( .A(n3989), .ZN(\xmem_inst/n3804 ) );
  OAI22_X1 U5324 ( .A1(n4004), .A2(s_data_in_x[19]), .B1(
        \xmem_inst/mem[42][19] ), .B2(n4003), .ZN(n3990) );
  INV_X1 U5325 ( .A(n3990), .ZN(\xmem_inst/n3805 ) );
  OAI22_X1 U5326 ( .A1(n4004), .A2(s_data_in_x[20]), .B1(
        \xmem_inst/mem[42][20] ), .B2(n4000), .ZN(n3991) );
  INV_X1 U5327 ( .A(n3991), .ZN(\xmem_inst/n3806 ) );
  OAI22_X1 U5328 ( .A1(n4004), .A2(s_data_in_x[21]), .B1(
        \xmem_inst/mem[42][21] ), .B2(n4000), .ZN(n3992) );
  INV_X1 U5329 ( .A(n3992), .ZN(\xmem_inst/n3807 ) );
  OAI22_X1 U5330 ( .A1(n4004), .A2(s_data_in_x[22]), .B1(
        \xmem_inst/mem[42][22] ), .B2(n4003), .ZN(n3993) );
  INV_X1 U5331 ( .A(n3993), .ZN(\xmem_inst/n3808 ) );
  OAI22_X1 U5332 ( .A1(n4004), .A2(s_data_in_x[23]), .B1(
        \xmem_inst/mem[42][23] ), .B2(n4003), .ZN(n3994) );
  INV_X1 U5333 ( .A(n3994), .ZN(\xmem_inst/n3809 ) );
  OAI22_X1 U5334 ( .A1(n4004), .A2(s_data_in_x[24]), .B1(
        \xmem_inst/mem[42][24] ), .B2(n4003), .ZN(n3995) );
  INV_X1 U5335 ( .A(n3995), .ZN(\xmem_inst/n3810 ) );
  OAI22_X1 U5336 ( .A1(n4004), .A2(s_data_in_x[25]), .B1(
        \xmem_inst/mem[42][25] ), .B2(n4000), .ZN(n3996) );
  INV_X1 U5337 ( .A(n3996), .ZN(\xmem_inst/n3811 ) );
  OAI22_X1 U5338 ( .A1(n4004), .A2(s_data_in_x[26]), .B1(
        \xmem_inst/mem[42][26] ), .B2(n4003), .ZN(n3997) );
  INV_X1 U5339 ( .A(n3997), .ZN(\xmem_inst/n3812 ) );
  OAI22_X1 U5340 ( .A1(n4004), .A2(s_data_in_x[27]), .B1(
        \xmem_inst/mem[42][27] ), .B2(n4000), .ZN(n3998) );
  INV_X1 U5341 ( .A(n3998), .ZN(\xmem_inst/n3813 ) );
  OAI22_X1 U5342 ( .A1(n4004), .A2(s_data_in_x[28]), .B1(
        \xmem_inst/mem[42][28] ), .B2(n4003), .ZN(n3999) );
  INV_X1 U5343 ( .A(n3999), .ZN(\xmem_inst/n3814 ) );
  OAI22_X1 U5344 ( .A1(n4004), .A2(s_data_in_x[29]), .B1(
        \xmem_inst/mem[42][29] ), .B2(n4000), .ZN(n4001) );
  INV_X1 U5345 ( .A(n4001), .ZN(\xmem_inst/n3815 ) );
  OAI22_X1 U5346 ( .A1(n4004), .A2(s_data_in_x[30]), .B1(
        \xmem_inst/mem[42][30] ), .B2(n4003), .ZN(n4002) );
  INV_X1 U5347 ( .A(n4002), .ZN(\xmem_inst/n3816 ) );
  OAI22_X1 U5348 ( .A1(n4004), .A2(s_data_in_x[31]), .B1(
        \xmem_inst/mem[42][31] ), .B2(n4003), .ZN(n4005) );
  INV_X1 U5349 ( .A(n4005), .ZN(\xmem_inst/n3817 ) );
  NAND4_X1 U5351 ( .A1(\ctrl_conv_output_inst/cnt_conv [2]), .A2(n4006), .A3(
        n4079), .A4(n4072), .ZN(n4008) );
  INV_X1 U5352 ( .A(reset), .ZN(n4023) );
  NAND4_X1 U5353 ( .A1(\ctrl_conv_output_inst/cnt_conv [4]), .A2(
        \ctrl_conv_output_inst/cnt_conv [3]), .A3(n4023), .A4(n4111), .ZN(
        n4007) );
  NOR2_X1 U5354 ( .A1(n4008), .A2(n4007), .ZN(\ctrl_conv_output_inst/N80 ) );
  NAND3_X1 U5355 ( .A1(n4009), .A2(n4023), .A3(n4010), .ZN(n4047) );
  INV_X1 U5356 ( .A(n4047), .ZN(\ctrl_conv_output_inst/N77 ) );
  NOR2_X1 U5357 ( .A1(s_ready_x), .A2(reset), .ZN(N23) );
  NAND2_X1 U5358 ( .A1(n4009), .A2(n4023), .ZN(n4046) );
  NAND3_X1 U5359 ( .A1(n4010), .A2(n4071), .A3(n4023), .ZN(n4011) );
  OAI22_X1 U5360 ( .A1(n4071), .A2(n4046), .B1(n4012), .B2(n4011), .ZN(n121)
         );
  OAI21_X1 U5361 ( .B1(\ctrl_conv_output_inst/m_pre_valid_y ), .B2(n4071), .A(
        n4025), .ZN(n4014) );
  AOI22_X1 U5362 ( .A1(\ctrl_conv_output_inst/cnt_conv [0]), .A2(n4014), .B1(
        n4013), .B2(n4072), .ZN(n119) );
  OAI21_X1 U5363 ( .B1(n4015), .B2(n4072), .A(n4025), .ZN(n4019) );
  NAND2_X1 U5364 ( .A1(n4016), .A2(n4079), .ZN(n4018) );
  OAI22_X1 U5365 ( .A1(n4019), .A2(n4079), .B1(n4072), .B2(n4018), .ZN(n118)
         );
  NAND4_X1 U5366 ( .A1(\ctrl_conv_output_inst/cnt_conv [1]), .A2(n4016), .A3(
        \ctrl_conv_output_inst/cnt_conv [0]), .A4(n4080), .ZN(n4017) );
  OAI221_X1 U5367 ( .B1(n4080), .B2(n4019), .C1(n4080), .C2(n4018), .A(n4017), 
        .ZN(n117) );
  INV_X1 U5368 ( .A(n4020), .ZN(n4022) );
  AOI22_X1 U5369 ( .A1(\ctrl_conv_output_inst/cnt_conv [4]), .A2(n4022), .B1(
        n4021), .B2(n4076), .ZN(n115) );
  NAND2_X1 U5370 ( .A1(m_valid_y), .A2(n4023), .ZN(n4024) );
  OAI22_X1 U5371 ( .A1(m_ready_y), .A2(n4024), .B1(n4047), .B2(n4075), .ZN(
        n114) );
  OAI21_X1 U5372 ( .B1(n4102), .B2(n4026), .A(n4025), .ZN(n113) );
  AOI22_X1 U5373 ( .A1(\ctrl_conv_output_inst/cnt_conv [0]), .A2(n4042), .B1(
        n4082), .B2(n4036), .ZN(n4027) );
  OAI21_X1 U5374 ( .B1(n4082), .B2(n4032), .A(n4027), .ZN(n112) );
  OR2_X1 U5375 ( .A1(xmem_addr[1]), .A2(n4041), .ZN(n4030) );
  OAI21_X1 U5376 ( .B1(xmem_addr[0]), .B2(n4041), .A(n4032), .ZN(n4028) );
  AOI22_X1 U5377 ( .A1(xmem_addr[1]), .A2(n4028), .B1(n4042), .B2(
        \ctrl_conv_output_inst/cnt_conv [1]), .ZN(n4029) );
  OAI21_X1 U5378 ( .B1(n4082), .B2(n4030), .A(n4029), .ZN(n111) );
  NAND4_X1 U5379 ( .A1(xmem_addr[2]), .A2(xmem_addr[0]), .A3(xmem_addr[1]), 
        .A4(n4036), .ZN(n4037) );
  NOR2_X1 U5380 ( .A1(n4105), .A2(n4031), .ZN(n4033) );
  OAI21_X1 U5381 ( .B1(n4041), .B2(n4033), .A(n4032), .ZN(n4035) );
  AOI22_X1 U5382 ( .A1(xmem_addr[3]), .A2(n4035), .B1(n4042), .B2(
        \ctrl_conv_output_inst/cnt_conv [3]), .ZN(n4034) );
  OAI21_X1 U5383 ( .B1(xmem_addr[3]), .B2(n4037), .A(n4034), .ZN(n109) );
  AOI21_X1 U5384 ( .B1(n4083), .B2(n4036), .A(n4035), .ZN(n4040) );
  NOR2_X1 U5385 ( .A1(n4083), .A2(n4037), .ZN(n4039) );
  AOI22_X1 U5386 ( .A1(\ctrl_conv_output_inst/cnt_conv [4]), .A2(n4042), .B1(
        n4039), .B2(n4081), .ZN(n4038) );
  OAI21_X1 U5387 ( .B1(n4040), .B2(n4081), .A(n4038), .ZN(n108) );
  NAND2_X1 U5388 ( .A1(n4039), .A2(xmem_addr[4]), .ZN(n4045) );
  OAI21_X1 U5389 ( .B1(xmem_addr[4]), .B2(n4041), .A(n4040), .ZN(n4043) );
  AOI22_X1 U5390 ( .A1(xmem_addr[5]), .A2(n4043), .B1(n4042), .B2(
        \ctrl_conv_output_inst/cnt_conv [5]), .ZN(n4044) );
  OAI21_X1 U5391 ( .B1(n4045), .B2(xmem_addr[5]), .A(n4044), .ZN(n107) );
  OAI22_X1 U5392 ( .A1(n4071), .A2(n4047), .B1(n4075), .B2(n4046), .ZN(n106)
         );
endmodule

