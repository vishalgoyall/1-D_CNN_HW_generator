
module conv_16_4_16_1 ( clk, reset, s_data_in_x, s_valid_x, s_ready_x, 
        m_data_out_y, m_valid_y, m_ready_y );
  input [15:0] s_data_in_x;
  output [15:0] m_data_out_y;
  input clk, reset, s_valid_x, m_ready_y;
  output s_ready_x, m_valid_y;
  wire   conv_done, N19, \xmem_inst/N29 , \xmem_inst/N28 , \xmem_inst/N27 ,
         \xmem_inst/N26 , \xmem_inst/N25 , \xmem_inst/N24 , \xmem_inst/N23 ,
         \xmem_inst/N22 , \xmem_inst/N21 , \xmem_inst/N20 , \xmem_inst/N19 ,
         \xmem_inst/N18 , \xmem_inst/N17 , \xmem_inst/N16 , \xmem_inst/N15 ,
         \xmem_inst/N14 , \xmem_inst/mem[15][15] , \xmem_inst/mem[15][14] ,
         \xmem_inst/mem[15][13] , \xmem_inst/mem[15][12] ,
         \xmem_inst/mem[15][11] , \xmem_inst/mem[15][10] ,
         \xmem_inst/mem[15][9] , \xmem_inst/mem[15][8] ,
         \xmem_inst/mem[15][7] , \xmem_inst/mem[15][6] ,
         \xmem_inst/mem[15][5] , \xmem_inst/mem[15][4] ,
         \xmem_inst/mem[15][3] , \xmem_inst/mem[15][2] ,
         \xmem_inst/mem[15][1] , \xmem_inst/mem[15][0] ,
         \xmem_inst/mem[14][15] , \xmem_inst/mem[14][14] ,
         \xmem_inst/mem[14][13] , \xmem_inst/mem[14][12] ,
         \xmem_inst/mem[14][11] , \xmem_inst/mem[14][10] ,
         \xmem_inst/mem[14][9] , \xmem_inst/mem[14][8] ,
         \xmem_inst/mem[14][7] , \xmem_inst/mem[14][6] ,
         \xmem_inst/mem[14][5] , \xmem_inst/mem[14][4] ,
         \xmem_inst/mem[14][3] , \xmem_inst/mem[14][2] ,
         \xmem_inst/mem[14][1] , \xmem_inst/mem[14][0] ,
         \xmem_inst/mem[13][15] , \xmem_inst/mem[13][14] ,
         \xmem_inst/mem[13][13] , \xmem_inst/mem[13][12] ,
         \xmem_inst/mem[13][11] , \xmem_inst/mem[13][10] ,
         \xmem_inst/mem[13][9] , \xmem_inst/mem[13][8] ,
         \xmem_inst/mem[13][7] , \xmem_inst/mem[13][6] ,
         \xmem_inst/mem[13][5] , \xmem_inst/mem[13][4] ,
         \xmem_inst/mem[13][3] , \xmem_inst/mem[13][2] ,
         \xmem_inst/mem[13][1] , \xmem_inst/mem[13][0] ,
         \xmem_inst/mem[12][15] , \xmem_inst/mem[12][14] ,
         \xmem_inst/mem[12][13] , \xmem_inst/mem[12][12] ,
         \xmem_inst/mem[12][11] , \xmem_inst/mem[12][10] ,
         \xmem_inst/mem[12][9] , \xmem_inst/mem[12][8] ,
         \xmem_inst/mem[12][7] , \xmem_inst/mem[12][6] ,
         \xmem_inst/mem[12][5] , \xmem_inst/mem[12][4] ,
         \xmem_inst/mem[12][3] , \xmem_inst/mem[12][2] ,
         \xmem_inst/mem[12][1] , \xmem_inst/mem[12][0] ,
         \xmem_inst/mem[11][15] , \xmem_inst/mem[11][14] ,
         \xmem_inst/mem[11][13] , \xmem_inst/mem[11][12] ,
         \xmem_inst/mem[11][11] , \xmem_inst/mem[11][10] ,
         \xmem_inst/mem[11][9] , \xmem_inst/mem[11][8] ,
         \xmem_inst/mem[11][7] , \xmem_inst/mem[11][6] ,
         \xmem_inst/mem[11][5] , \xmem_inst/mem[11][4] ,
         \xmem_inst/mem[11][3] , \xmem_inst/mem[11][2] ,
         \xmem_inst/mem[11][1] , \xmem_inst/mem[11][0] ,
         \xmem_inst/mem[10][15] , \xmem_inst/mem[10][14] ,
         \xmem_inst/mem[10][13] , \xmem_inst/mem[10][12] ,
         \xmem_inst/mem[10][11] , \xmem_inst/mem[10][10] ,
         \xmem_inst/mem[10][9] , \xmem_inst/mem[10][8] ,
         \xmem_inst/mem[10][7] , \xmem_inst/mem[10][6] ,
         \xmem_inst/mem[10][5] , \xmem_inst/mem[10][4] ,
         \xmem_inst/mem[10][3] , \xmem_inst/mem[10][2] ,
         \xmem_inst/mem[10][1] , \xmem_inst/mem[10][0] ,
         \xmem_inst/mem[9][15] , \xmem_inst/mem[9][14] ,
         \xmem_inst/mem[9][13] , \xmem_inst/mem[9][12] ,
         \xmem_inst/mem[9][11] , \xmem_inst/mem[9][10] , \xmem_inst/mem[9][9] ,
         \xmem_inst/mem[9][8] , \xmem_inst/mem[9][7] , \xmem_inst/mem[9][6] ,
         \xmem_inst/mem[9][5] , \xmem_inst/mem[9][4] , \xmem_inst/mem[9][3] ,
         \xmem_inst/mem[9][2] , \xmem_inst/mem[9][1] , \xmem_inst/mem[9][0] ,
         \xmem_inst/mem[8][15] , \xmem_inst/mem[8][14] ,
         \xmem_inst/mem[8][13] , \xmem_inst/mem[8][12] ,
         \xmem_inst/mem[8][11] , \xmem_inst/mem[8][10] , \xmem_inst/mem[8][9] ,
         \xmem_inst/mem[8][8] , \xmem_inst/mem[8][7] , \xmem_inst/mem[8][6] ,
         \xmem_inst/mem[8][5] , \xmem_inst/mem[8][4] , \xmem_inst/mem[8][3] ,
         \xmem_inst/mem[8][2] , \xmem_inst/mem[8][1] , \xmem_inst/mem[8][0] ,
         \xmem_inst/mem[6][15] , \xmem_inst/mem[6][14] ,
         \xmem_inst/mem[6][13] , \xmem_inst/mem[6][12] ,
         \xmem_inst/mem[6][11] , \xmem_inst/mem[6][10] , \xmem_inst/mem[6][9] ,
         \xmem_inst/mem[6][8] , \xmem_inst/mem[6][7] , \xmem_inst/mem[6][6] ,
         \xmem_inst/mem[6][5] , \xmem_inst/mem[6][4] , \xmem_inst/mem[6][3] ,
         \xmem_inst/mem[6][2] , \xmem_inst/mem[6][1] , \xmem_inst/mem[6][0] ,
         \xmem_inst/mem[5][15] , \xmem_inst/mem[5][14] ,
         \xmem_inst/mem[5][13] , \xmem_inst/mem[5][12] ,
         \xmem_inst/mem[5][11] , \xmem_inst/mem[5][10] , \xmem_inst/mem[5][9] ,
         \xmem_inst/mem[5][8] , \xmem_inst/mem[5][7] , \xmem_inst/mem[5][6] ,
         \xmem_inst/mem[5][5] , \xmem_inst/mem[5][4] , \xmem_inst/mem[5][3] ,
         \xmem_inst/mem[5][2] , \xmem_inst/mem[5][1] , \xmem_inst/mem[5][0] ,
         \xmem_inst/mem[4][15] , \xmem_inst/mem[4][14] ,
         \xmem_inst/mem[4][13] , \xmem_inst/mem[4][12] ,
         \xmem_inst/mem[4][11] , \xmem_inst/mem[4][10] , \xmem_inst/mem[4][9] ,
         \xmem_inst/mem[4][8] , \xmem_inst/mem[4][7] , \xmem_inst/mem[4][6] ,
         \xmem_inst/mem[4][5] , \xmem_inst/mem[4][4] , \xmem_inst/mem[4][3] ,
         \xmem_inst/mem[4][2] , \xmem_inst/mem[4][1] , \xmem_inst/mem[4][0] ,
         \xmem_inst/mem[3][15] , \xmem_inst/mem[3][14] ,
         \xmem_inst/mem[3][13] , \xmem_inst/mem[3][12] ,
         \xmem_inst/mem[3][11] , \xmem_inst/mem[3][10] , \xmem_inst/mem[3][9] ,
         \xmem_inst/mem[3][8] , \xmem_inst/mem[3][7] , \xmem_inst/mem[3][6] ,
         \xmem_inst/mem[3][5] , \xmem_inst/mem[3][4] , \xmem_inst/mem[3][3] ,
         \xmem_inst/mem[3][2] , \xmem_inst/mem[3][1] , \xmem_inst/mem[3][0] ,
         \xmem_inst/mem[2][15] , \xmem_inst/mem[2][14] ,
         \xmem_inst/mem[2][13] , \xmem_inst/mem[2][12] ,
         \xmem_inst/mem[2][11] , \xmem_inst/mem[2][10] , \xmem_inst/mem[2][9] ,
         \xmem_inst/mem[2][8] , \xmem_inst/mem[2][7] , \xmem_inst/mem[2][6] ,
         \xmem_inst/mem[2][5] , \xmem_inst/mem[2][4] , \xmem_inst/mem[2][3] ,
         \xmem_inst/mem[2][2] , \xmem_inst/mem[2][1] , \xmem_inst/mem[2][0] ,
         \xmem_inst/mem[1][15] , \xmem_inst/mem[1][14] ,
         \xmem_inst/mem[1][13] , \xmem_inst/mem[1][12] ,
         \xmem_inst/mem[1][11] , \xmem_inst/mem[1][10] , \xmem_inst/mem[1][9] ,
         \xmem_inst/mem[1][8] , \xmem_inst/mem[1][7] , \xmem_inst/mem[1][6] ,
         \xmem_inst/mem[1][5] , \xmem_inst/mem[1][4] , \xmem_inst/mem[1][3] ,
         \xmem_inst/mem[1][2] , \xmem_inst/mem[1][1] , \xmem_inst/mem[1][0] ,
         \xmem_inst/mem[0][15] , \xmem_inst/mem[0][14] ,
         \xmem_inst/mem[0][13] , \xmem_inst/mem[0][12] ,
         \xmem_inst/mem[0][11] , \xmem_inst/mem[0][10] , \xmem_inst/mem[0][9] ,
         \xmem_inst/mem[0][8] , \xmem_inst/mem[0][7] , \xmem_inst/mem[0][6] ,
         \xmem_inst/mem[0][5] , \xmem_inst/mem[0][4] , \xmem_inst/mem[0][3] ,
         \xmem_inst/mem[0][2] , \xmem_inst/mem[0][1] , \xmem_inst/mem[0][0] ,
         \fmem_inst/N14 , \fmem_inst/N13 , \fmem_inst/N12 ,
         \ctrl_conv_output_inst/N74 , \ctrl_conv_output_inst/m_pre_valid_y ,
         \ctrl_conv_output_inst/conv_start_accum ,
         \ctrl_conv_output_inst/m_pre_pre_valid_y , n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133;
  wire   [3:0] xmem_addr;
  wire   [15:0] xmem_data;
  wire   [15:0] fmem_data;
  wire   [3:0] \ctrl_conv_output_inst/cnt_conv ;
  wire   [15:0] \mac_unit_inst/adder_reg ;
  wire   [15:0] \mac_unit_inst/x_mult_f_reg ;
  assign m_data_out_y[15] = 1'b0;

  DFF_X1 \xmem_inst/data_out_reg[2]  ( .D(\xmem_inst/N27 ), .CK(clk), .QN(
        n1831) );
  DFF_X1 \xmem_inst/data_out_reg[3]  ( .D(\xmem_inst/N26 ), .CK(clk), .QN(
        n1832) );
  DFF_X1 \xmem_inst/data_out_reg[6]  ( .D(\xmem_inst/N23 ), .CK(clk), .Q(
        xmem_data[6]), .QN(n911) );
  DFF_X1 \xmem_inst/data_out_reg[7]  ( .D(\xmem_inst/N22 ), .CK(clk), .Q(
        xmem_data[7]), .QN(n908) );
  DFF_X1 \xmem_inst/data_out_reg[8]  ( .D(\xmem_inst/N21 ), .CK(clk), .QN(
        n1815) );
  DFF_X1 \xmem_inst/data_out_reg[9]  ( .D(\xmem_inst/N20 ), .CK(clk), .Q(
        xmem_data[9]), .QN(n909) );
  DFF_X1 \xmem_inst/data_out_reg[10]  ( .D(\xmem_inst/N19 ), .CK(clk), .Q(
        xmem_data[10]), .QN(n1818) );
  DFF_X1 \xmem_inst/data_out_reg[12]  ( .D(\xmem_inst/N17 ), .CK(clk), .Q(
        xmem_data[12]), .QN(n906) );
  DFF_X1 \xmem_inst/data_out_reg[13]  ( .D(\xmem_inst/N16 ), .CK(clk), .Q(
        xmem_data[13]), .QN(n1817) );
  DFF_X1 \xmem_inst/data_out_reg[14]  ( .D(\xmem_inst/N15 ), .CK(clk), .Q(
        xmem_data[14]), .QN(n907) );
  DFF_X1 \fmem_inst/z_reg[4]  ( .D(\fmem_inst/N14 ), .CK(clk), .Q(fmem_data[4]), .QN(n1820) );
  DFF_X1 \fmem_inst/z_reg[15]  ( .D(n1834), .CK(clk), .Q(fmem_data[15]), .QN(
        n1819) );
  DFF_X1 \ctrl_conv_output_inst/conv_done_reg  ( .D(
        \ctrl_conv_output_inst/N74 ), .CK(clk), .Q(conv_done) );
  DFF_X1 \ctrl_conv_output_inst/m_pre_pre_valid_y_reg  ( .D(n879), .CK(clk), 
        .Q(\ctrl_conv_output_inst/m_pre_pre_valid_y ), .QN(n1836) );
  DFF_X1 \ctrl_conv_output_inst/m_pre_valid_y_reg  ( .D(n612), .CK(clk), .Q(
        \ctrl_conv_output_inst/m_pre_valid_y ), .QN(n1870) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[0]  ( .D(n877), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [0]), .QN(n1841) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[1]  ( .D(n876), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [1]), .QN(n1840) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[2]  ( .D(n875), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [2]), .QN(n1837) );
  DFF_X1 \ctrl_conv_output_inst/m_valid_y_reg  ( .D(n874), .CK(clk), .Q(
        m_valid_y), .QN(n2035) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[3]  ( .D(n869), .CK(clk), .Q(
        xmem_addr[3]), .QN(n1842) );
  DFF_X1 \ctrl_xmem_write_inst/s_ready_reg  ( .D(n873), .CK(clk), .Q(s_ready_x), .QN(n2116) );
  DFF_X1 conv_pre_start_reg ( .D(N19), .CK(clk), .QN(n2117) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[0]  ( .D(n872), .CK(clk), .Q(
        xmem_addr[0]), .QN(n1833) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[1]  ( .D(n871), .CK(clk), .Q(
        xmem_addr[1]), .QN(n1838) );
  DFF_X1 \xmem_inst/mem_reg[12][0]  ( .D(n676), .CK(clk), .Q(
        \xmem_inst/mem[12][0] ), .QN(n2084) );
  DFF_X1 \xmem_inst/mem_reg[12][1]  ( .D(n675), .CK(clk), .Q(
        \xmem_inst/mem[12][1] ), .QN(n2085) );
  DFF_X1 \xmem_inst/mem_reg[12][2]  ( .D(n674), .CK(clk), .Q(
        \xmem_inst/mem[12][2] ), .QN(n2086) );
  DFF_X1 \xmem_inst/mem_reg[12][3]  ( .D(n673), .CK(clk), .Q(
        \xmem_inst/mem[12][3] ), .QN(n2087) );
  DFF_X1 \xmem_inst/mem_reg[12][4]  ( .D(n672), .CK(clk), .Q(
        \xmem_inst/mem[12][4] ), .QN(n2088) );
  DFF_X1 \xmem_inst/mem_reg[12][5]  ( .D(n671), .CK(clk), .Q(
        \xmem_inst/mem[12][5] ), .QN(n2089) );
  DFF_X1 \xmem_inst/mem_reg[12][6]  ( .D(n670), .CK(clk), .Q(
        \xmem_inst/mem[12][6] ), .QN(n2090) );
  DFF_X1 \xmem_inst/mem_reg[12][7]  ( .D(n669), .CK(clk), .Q(
        \xmem_inst/mem[12][7] ), .QN(n2091) );
  DFF_X1 \xmem_inst/mem_reg[12][8]  ( .D(n668), .CK(clk), .Q(
        \xmem_inst/mem[12][8] ), .QN(n2092) );
  DFF_X1 \xmem_inst/mem_reg[12][9]  ( .D(n667), .CK(clk), .Q(
        \xmem_inst/mem[12][9] ), .QN(n2093) );
  DFF_X1 \xmem_inst/mem_reg[12][10]  ( .D(n666), .CK(clk), .Q(
        \xmem_inst/mem[12][10] ), .QN(n2094) );
  DFF_X1 \xmem_inst/mem_reg[12][11]  ( .D(n665), .CK(clk), .Q(
        \xmem_inst/mem[12][11] ), .QN(n2095) );
  DFF_X1 \xmem_inst/mem_reg[12][12]  ( .D(n664), .CK(clk), .Q(
        \xmem_inst/mem[12][12] ), .QN(n2096) );
  DFF_X1 \xmem_inst/mem_reg[12][13]  ( .D(n663), .CK(clk), .Q(
        \xmem_inst/mem[12][13] ), .QN(n2097) );
  DFF_X1 \xmem_inst/mem_reg[12][14]  ( .D(n662), .CK(clk), .Q(
        \xmem_inst/mem[12][14] ), .QN(n2098) );
  DFF_X1 \xmem_inst/mem_reg[12][15]  ( .D(n661), .CK(clk), .Q(
        \xmem_inst/mem[12][15] ), .QN(n2099) );
  DFF_X1 \xmem_inst/mem_reg[13][0]  ( .D(n660), .CK(clk), .Q(
        \xmem_inst/mem[13][0] ), .QN(n2003) );
  DFF_X1 \xmem_inst/mem_reg[13][1]  ( .D(n659), .CK(clk), .Q(
        \xmem_inst/mem[13][1] ), .QN(n2004) );
  DFF_X1 \xmem_inst/mem_reg[13][2]  ( .D(n658), .CK(clk), .Q(
        \xmem_inst/mem[13][2] ), .QN(n2005) );
  DFF_X1 \xmem_inst/mem_reg[13][3]  ( .D(n657), .CK(clk), .Q(
        \xmem_inst/mem[13][3] ), .QN(n2006) );
  DFF_X1 \xmem_inst/mem_reg[13][4]  ( .D(n656), .CK(clk), .Q(
        \xmem_inst/mem[13][4] ), .QN(n2007) );
  DFF_X1 \xmem_inst/mem_reg[13][5]  ( .D(n655), .CK(clk), .Q(
        \xmem_inst/mem[13][5] ), .QN(n2008) );
  DFF_X1 \xmem_inst/mem_reg[13][6]  ( .D(n654), .CK(clk), .Q(
        \xmem_inst/mem[13][6] ), .QN(n2009) );
  DFF_X1 \xmem_inst/mem_reg[13][7]  ( .D(n653), .CK(clk), .Q(
        \xmem_inst/mem[13][7] ), .QN(n2010) );
  DFF_X1 \xmem_inst/mem_reg[13][8]  ( .D(n652), .CK(clk), .Q(
        \xmem_inst/mem[13][8] ), .QN(n2011) );
  DFF_X1 \xmem_inst/mem_reg[13][9]  ( .D(n651), .CK(clk), .Q(
        \xmem_inst/mem[13][9] ), .QN(n2012) );
  DFF_X1 \xmem_inst/mem_reg[13][10]  ( .D(n650), .CK(clk), .Q(
        \xmem_inst/mem[13][10] ), .QN(n2013) );
  DFF_X1 \xmem_inst/mem_reg[13][11]  ( .D(n649), .CK(clk), .Q(
        \xmem_inst/mem[13][11] ), .QN(n2014) );
  DFF_X1 \xmem_inst/mem_reg[13][12]  ( .D(n648), .CK(clk), .Q(
        \xmem_inst/mem[13][12] ), .QN(n2015) );
  DFF_X1 \xmem_inst/mem_reg[13][13]  ( .D(n647), .CK(clk), .Q(
        \xmem_inst/mem[13][13] ), .QN(n2016) );
  DFF_X1 \xmem_inst/mem_reg[13][14]  ( .D(n646), .CK(clk), .Q(
        \xmem_inst/mem[13][14] ), .QN(n2017) );
  DFF_X1 \xmem_inst/mem_reg[13][15]  ( .D(n645), .CK(clk), .Q(
        \xmem_inst/mem[13][15] ), .QN(n2018) );
  DFF_X1 \xmem_inst/mem_reg[14][0]  ( .D(n644), .CK(clk), .Q(
        \xmem_inst/mem[14][0] ), .QN(n2100) );
  DFF_X1 \xmem_inst/mem_reg[14][1]  ( .D(n643), .CK(clk), .Q(
        \xmem_inst/mem[14][1] ), .QN(n2101) );
  DFF_X1 \xmem_inst/mem_reg[14][2]  ( .D(n642), .CK(clk), .Q(
        \xmem_inst/mem[14][2] ), .QN(n2102) );
  DFF_X1 \xmem_inst/mem_reg[14][3]  ( .D(n641), .CK(clk), .Q(
        \xmem_inst/mem[14][3] ), .QN(n2103) );
  DFF_X1 \xmem_inst/mem_reg[14][4]  ( .D(n640), .CK(clk), .Q(
        \xmem_inst/mem[14][4] ), .QN(n2104) );
  DFF_X1 \xmem_inst/mem_reg[14][5]  ( .D(n639), .CK(clk), .Q(
        \xmem_inst/mem[14][5] ), .QN(n2105) );
  DFF_X1 \xmem_inst/mem_reg[14][6]  ( .D(n638), .CK(clk), .Q(
        \xmem_inst/mem[14][6] ), .QN(n2106) );
  DFF_X1 \xmem_inst/mem_reg[14][7]  ( .D(n637), .CK(clk), .Q(
        \xmem_inst/mem[14][7] ), .QN(n2107) );
  DFF_X1 \xmem_inst/mem_reg[14][8]  ( .D(n636), .CK(clk), .Q(
        \xmem_inst/mem[14][8] ), .QN(n2108) );
  DFF_X1 \xmem_inst/mem_reg[14][9]  ( .D(n635), .CK(clk), .Q(
        \xmem_inst/mem[14][9] ), .QN(n2109) );
  DFF_X1 \xmem_inst/mem_reg[14][10]  ( .D(n634), .CK(clk), .Q(
        \xmem_inst/mem[14][10] ), .QN(n2110) );
  DFF_X1 \xmem_inst/mem_reg[14][11]  ( .D(n633), .CK(clk), .Q(
        \xmem_inst/mem[14][11] ), .QN(n2111) );
  DFF_X1 \xmem_inst/mem_reg[14][12]  ( .D(n632), .CK(clk), .Q(
        \xmem_inst/mem[14][12] ), .QN(n2112) );
  DFF_X1 \xmem_inst/mem_reg[14][13]  ( .D(n631), .CK(clk), .Q(
        \xmem_inst/mem[14][13] ), .QN(n2113) );
  DFF_X1 \xmem_inst/mem_reg[14][14]  ( .D(n630), .CK(clk), .Q(
        \xmem_inst/mem[14][14] ), .QN(n2114) );
  DFF_X1 \xmem_inst/mem_reg[14][15]  ( .D(n629), .CK(clk), .Q(
        \xmem_inst/mem[14][15] ), .QN(n2115) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[2]  ( .D(n870), .CK(clk), .Q(
        xmem_addr[2]), .QN(n1835) );
  DFF_X1 \xmem_inst/mem_reg[4][0]  ( .D(n804), .CK(clk), .Q(
        \xmem_inst/mem[4][0] ), .QN(n2068) );
  DFF_X1 \xmem_inst/mem_reg[4][1]  ( .D(n803), .CK(clk), .Q(
        \xmem_inst/mem[4][1] ), .QN(n2069) );
  DFF_X1 \xmem_inst/mem_reg[4][2]  ( .D(n802), .CK(clk), .Q(
        \xmem_inst/mem[4][2] ), .QN(n2070) );
  DFF_X1 \xmem_inst/mem_reg[4][3]  ( .D(n801), .CK(clk), .Q(
        \xmem_inst/mem[4][3] ), .QN(n2071) );
  DFF_X1 \xmem_inst/mem_reg[4][4]  ( .D(n800), .CK(clk), .Q(
        \xmem_inst/mem[4][4] ), .QN(n2072) );
  DFF_X1 \xmem_inst/mem_reg[4][5]  ( .D(n799), .CK(clk), .Q(
        \xmem_inst/mem[4][5] ), .QN(n2073) );
  DFF_X1 \xmem_inst/mem_reg[4][6]  ( .D(n798), .CK(clk), .Q(
        \xmem_inst/mem[4][6] ), .QN(n2074) );
  DFF_X1 \xmem_inst/mem_reg[4][7]  ( .D(n797), .CK(clk), .Q(
        \xmem_inst/mem[4][7] ), .QN(n2075) );
  DFF_X1 \xmem_inst/mem_reg[4][8]  ( .D(n796), .CK(clk), .Q(
        \xmem_inst/mem[4][8] ), .QN(n2076) );
  DFF_X1 \xmem_inst/mem_reg[4][9]  ( .D(n795), .CK(clk), .Q(
        \xmem_inst/mem[4][9] ), .QN(n2077) );
  DFF_X1 \xmem_inst/mem_reg[4][10]  ( .D(n794), .CK(clk), .Q(
        \xmem_inst/mem[4][10] ), .QN(n2078) );
  DFF_X1 \xmem_inst/mem_reg[4][11]  ( .D(n793), .CK(clk), .Q(
        \xmem_inst/mem[4][11] ), .QN(n2079) );
  DFF_X1 \xmem_inst/mem_reg[4][12]  ( .D(n792), .CK(clk), .Q(
        \xmem_inst/mem[4][12] ), .QN(n2080) );
  DFF_X1 \xmem_inst/mem_reg[4][13]  ( .D(n791), .CK(clk), .Q(
        \xmem_inst/mem[4][13] ), .QN(n2081) );
  DFF_X1 \xmem_inst/mem_reg[4][14]  ( .D(n790), .CK(clk), .Q(
        \xmem_inst/mem[4][14] ), .QN(n2082) );
  DFF_X1 \xmem_inst/mem_reg[4][15]  ( .D(n789), .CK(clk), .Q(
        \xmem_inst/mem[4][15] ), .QN(n2083) );
  DFF_X1 \xmem_inst/mem_reg[5][0]  ( .D(n788), .CK(clk), .Q(
        \xmem_inst/mem[5][0] ), .QN(n1987) );
  DFF_X1 \xmem_inst/mem_reg[5][1]  ( .D(n787), .CK(clk), .Q(
        \xmem_inst/mem[5][1] ), .QN(n1988) );
  DFF_X1 \xmem_inst/mem_reg[5][2]  ( .D(n786), .CK(clk), .Q(
        \xmem_inst/mem[5][2] ), .QN(n1989) );
  DFF_X1 \xmem_inst/mem_reg[5][3]  ( .D(n785), .CK(clk), .Q(
        \xmem_inst/mem[5][3] ), .QN(n1990) );
  DFF_X1 \xmem_inst/mem_reg[5][4]  ( .D(n784), .CK(clk), .Q(
        \xmem_inst/mem[5][4] ), .QN(n1991) );
  DFF_X1 \xmem_inst/mem_reg[5][5]  ( .D(n783), .CK(clk), .Q(
        \xmem_inst/mem[5][5] ), .QN(n1992) );
  DFF_X1 \xmem_inst/mem_reg[5][6]  ( .D(n782), .CK(clk), .Q(
        \xmem_inst/mem[5][6] ), .QN(n1993) );
  DFF_X1 \xmem_inst/mem_reg[5][7]  ( .D(n781), .CK(clk), .Q(
        \xmem_inst/mem[5][7] ), .QN(n1994) );
  DFF_X1 \xmem_inst/mem_reg[5][8]  ( .D(n780), .CK(clk), .Q(
        \xmem_inst/mem[5][8] ), .QN(n1995) );
  DFF_X1 \xmem_inst/mem_reg[5][9]  ( .D(n779), .CK(clk), .Q(
        \xmem_inst/mem[5][9] ), .QN(n1996) );
  DFF_X1 \xmem_inst/mem_reg[5][10]  ( .D(n778), .CK(clk), .Q(
        \xmem_inst/mem[5][10] ), .QN(n1997) );
  DFF_X1 \xmem_inst/mem_reg[5][11]  ( .D(n777), .CK(clk), .Q(
        \xmem_inst/mem[5][11] ), .QN(n1998) );
  DFF_X1 \xmem_inst/mem_reg[5][12]  ( .D(n776), .CK(clk), .Q(
        \xmem_inst/mem[5][12] ), .QN(n1999) );
  DFF_X1 \xmem_inst/mem_reg[5][13]  ( .D(n775), .CK(clk), .Q(
        \xmem_inst/mem[5][13] ), .QN(n2000) );
  DFF_X1 \xmem_inst/mem_reg[5][14]  ( .D(n774), .CK(clk), .Q(
        \xmem_inst/mem[5][14] ), .QN(n2001) );
  DFF_X1 \xmem_inst/mem_reg[5][15]  ( .D(n773), .CK(clk), .Q(
        \xmem_inst/mem[5][15] ), .QN(n2002) );
  DFF_X1 \xmem_inst/mem_reg[6][0]  ( .D(n772), .CK(clk), .Q(
        \xmem_inst/mem[6][0] ), .QN(n1939) );
  DFF_X1 \xmem_inst/mem_reg[6][1]  ( .D(n771), .CK(clk), .Q(
        \xmem_inst/mem[6][1] ), .QN(n1940) );
  DFF_X1 \xmem_inst/mem_reg[6][2]  ( .D(n770), .CK(clk), .Q(
        \xmem_inst/mem[6][2] ), .QN(n1941) );
  DFF_X1 \xmem_inst/mem_reg[6][3]  ( .D(n769), .CK(clk), .Q(
        \xmem_inst/mem[6][3] ), .QN(n1942) );
  DFF_X1 \xmem_inst/mem_reg[6][4]  ( .D(n768), .CK(clk), .Q(
        \xmem_inst/mem[6][4] ), .QN(n1943) );
  DFF_X1 \xmem_inst/mem_reg[6][5]  ( .D(n767), .CK(clk), .Q(
        \xmem_inst/mem[6][5] ), .QN(n1944) );
  DFF_X1 \xmem_inst/mem_reg[6][6]  ( .D(n766), .CK(clk), .Q(
        \xmem_inst/mem[6][6] ), .QN(n1945) );
  DFF_X1 \xmem_inst/mem_reg[6][7]  ( .D(n765), .CK(clk), .Q(
        \xmem_inst/mem[6][7] ), .QN(n1946) );
  DFF_X1 \xmem_inst/mem_reg[6][8]  ( .D(n764), .CK(clk), .Q(
        \xmem_inst/mem[6][8] ), .QN(n1947) );
  DFF_X1 \xmem_inst/mem_reg[6][9]  ( .D(n763), .CK(clk), .Q(
        \xmem_inst/mem[6][9] ), .QN(n1948) );
  DFF_X1 \xmem_inst/mem_reg[6][10]  ( .D(n762), .CK(clk), .Q(
        \xmem_inst/mem[6][10] ), .QN(n1949) );
  DFF_X1 \xmem_inst/mem_reg[6][11]  ( .D(n761), .CK(clk), .Q(
        \xmem_inst/mem[6][11] ), .QN(n1950) );
  DFF_X1 \xmem_inst/mem_reg[6][12]  ( .D(n760), .CK(clk), .Q(
        \xmem_inst/mem[6][12] ), .QN(n1951) );
  DFF_X1 \xmem_inst/mem_reg[6][13]  ( .D(n759), .CK(clk), .Q(
        \xmem_inst/mem[6][13] ), .QN(n1952) );
  DFF_X1 \xmem_inst/mem_reg[6][14]  ( .D(n758), .CK(clk), .Q(
        \xmem_inst/mem[6][14] ), .QN(n1953) );
  DFF_X1 \xmem_inst/mem_reg[6][15]  ( .D(n757), .CK(clk), .Q(
        \xmem_inst/mem[6][15] ), .QN(n1954) );
  DFF_X1 \xmem_inst/mem_reg[7][0]  ( .D(n756), .CK(clk), .QN(n1848) );
  DFF_X1 \xmem_inst/mem_reg[7][1]  ( .D(n755), .CK(clk), .QN(n1849) );
  DFF_X1 \xmem_inst/mem_reg[7][2]  ( .D(n754), .CK(clk), .QN(n1850) );
  DFF_X1 \xmem_inst/mem_reg[7][3]  ( .D(n753), .CK(clk), .QN(n1851) );
  DFF_X1 \xmem_inst/mem_reg[7][4]  ( .D(n752), .CK(clk), .QN(n1852) );
  DFF_X1 \xmem_inst/mem_reg[7][5]  ( .D(n751), .CK(clk), .QN(n1853) );
  DFF_X1 \xmem_inst/mem_reg[7][6]  ( .D(n750), .CK(clk), .QN(n1854) );
  DFF_X1 \xmem_inst/mem_reg[7][7]  ( .D(n749), .CK(clk), .QN(n1855) );
  DFF_X1 \xmem_inst/mem_reg[7][8]  ( .D(n748), .CK(clk), .QN(n1856) );
  DFF_X1 \xmem_inst/mem_reg[7][9]  ( .D(n747), .CK(clk), .QN(n1857) );
  DFF_X1 \xmem_inst/mem_reg[7][10]  ( .D(n746), .CK(clk), .QN(n1858) );
  DFF_X1 \xmem_inst/mem_reg[7][11]  ( .D(n745), .CK(clk), .QN(n1859) );
  DFF_X1 \xmem_inst/mem_reg[7][12]  ( .D(n744), .CK(clk), .QN(n1860) );
  DFF_X1 \xmem_inst/mem_reg[7][13]  ( .D(n743), .CK(clk), .QN(n1861) );
  DFF_X1 \xmem_inst/mem_reg[7][14]  ( .D(n742), .CK(clk), .QN(n1862) );
  DFF_X1 \xmem_inst/mem_reg[7][15]  ( .D(n741), .CK(clk), .QN(n1863) );
  DFF_X1 \xmem_inst/mem_reg[0][0]  ( .D(n868), .CK(clk), .Q(
        \xmem_inst/mem[0][0] ), .QN(n2036) );
  DFF_X1 \xmem_inst/mem_reg[0][1]  ( .D(n867), .CK(clk), .Q(
        \xmem_inst/mem[0][1] ), .QN(n2037) );
  DFF_X1 \xmem_inst/mem_reg[0][2]  ( .D(n866), .CK(clk), .Q(
        \xmem_inst/mem[0][2] ), .QN(n2038) );
  DFF_X1 \xmem_inst/mem_reg[0][3]  ( .D(n865), .CK(clk), .Q(
        \xmem_inst/mem[0][3] ), .QN(n2039) );
  DFF_X1 \xmem_inst/mem_reg[0][4]  ( .D(n864), .CK(clk), .Q(
        \xmem_inst/mem[0][4] ), .QN(n2040) );
  DFF_X1 \xmem_inst/mem_reg[0][5]  ( .D(n863), .CK(clk), .Q(
        \xmem_inst/mem[0][5] ), .QN(n2041) );
  DFF_X1 \xmem_inst/mem_reg[0][6]  ( .D(n862), .CK(clk), .Q(
        \xmem_inst/mem[0][6] ), .QN(n2042) );
  DFF_X1 \xmem_inst/mem_reg[0][7]  ( .D(n861), .CK(clk), .Q(
        \xmem_inst/mem[0][7] ), .QN(n2043) );
  DFF_X1 \xmem_inst/mem_reg[0][8]  ( .D(n860), .CK(clk), .Q(
        \xmem_inst/mem[0][8] ), .QN(n2044) );
  DFF_X1 \xmem_inst/mem_reg[0][9]  ( .D(n859), .CK(clk), .Q(
        \xmem_inst/mem[0][9] ), .QN(n2045) );
  DFF_X1 \xmem_inst/mem_reg[0][10]  ( .D(n858), .CK(clk), .Q(
        \xmem_inst/mem[0][10] ), .QN(n2046) );
  DFF_X1 \xmem_inst/mem_reg[0][11]  ( .D(n857), .CK(clk), .Q(
        \xmem_inst/mem[0][11] ), .QN(n2047) );
  DFF_X1 \xmem_inst/mem_reg[0][12]  ( .D(n856), .CK(clk), .Q(
        \xmem_inst/mem[0][12] ), .QN(n2048) );
  DFF_X1 \xmem_inst/mem_reg[0][13]  ( .D(n855), .CK(clk), .Q(
        \xmem_inst/mem[0][13] ), .QN(n2049) );
  DFF_X1 \xmem_inst/mem_reg[0][14]  ( .D(n854), .CK(clk), .Q(
        \xmem_inst/mem[0][14] ), .QN(n2050) );
  DFF_X1 \xmem_inst/mem_reg[0][15]  ( .D(n853), .CK(clk), .Q(
        \xmem_inst/mem[0][15] ), .QN(n2051) );
  DFF_X1 \xmem_inst/mem_reg[1][0]  ( .D(n852), .CK(clk), .Q(
        \xmem_inst/mem[1][0] ), .QN(n1955) );
  DFF_X1 \xmem_inst/mem_reg[1][1]  ( .D(n851), .CK(clk), .Q(
        \xmem_inst/mem[1][1] ), .QN(n1956) );
  DFF_X1 \xmem_inst/mem_reg[1][2]  ( .D(n850), .CK(clk), .Q(
        \xmem_inst/mem[1][2] ), .QN(n1957) );
  DFF_X1 \xmem_inst/mem_reg[1][3]  ( .D(n849), .CK(clk), .Q(
        \xmem_inst/mem[1][3] ), .QN(n1958) );
  DFF_X1 \xmem_inst/mem_reg[1][4]  ( .D(n848), .CK(clk), .Q(
        \xmem_inst/mem[1][4] ), .QN(n1959) );
  DFF_X1 \xmem_inst/mem_reg[1][5]  ( .D(n847), .CK(clk), .Q(
        \xmem_inst/mem[1][5] ), .QN(n1960) );
  DFF_X1 \xmem_inst/mem_reg[1][6]  ( .D(n846), .CK(clk), .Q(
        \xmem_inst/mem[1][6] ), .QN(n1961) );
  DFF_X1 \xmem_inst/mem_reg[1][7]  ( .D(n845), .CK(clk), .Q(
        \xmem_inst/mem[1][7] ), .QN(n1962) );
  DFF_X1 \xmem_inst/mem_reg[1][8]  ( .D(n844), .CK(clk), .Q(
        \xmem_inst/mem[1][8] ), .QN(n1963) );
  DFF_X1 \xmem_inst/mem_reg[1][9]  ( .D(n843), .CK(clk), .Q(
        \xmem_inst/mem[1][9] ), .QN(n1964) );
  DFF_X1 \xmem_inst/mem_reg[1][10]  ( .D(n842), .CK(clk), .Q(
        \xmem_inst/mem[1][10] ), .QN(n1965) );
  DFF_X1 \xmem_inst/mem_reg[1][11]  ( .D(n841), .CK(clk), .Q(
        \xmem_inst/mem[1][11] ), .QN(n1966) );
  DFF_X1 \xmem_inst/mem_reg[1][12]  ( .D(n840), .CK(clk), .Q(
        \xmem_inst/mem[1][12] ), .QN(n1967) );
  DFF_X1 \xmem_inst/mem_reg[1][13]  ( .D(n839), .CK(clk), .Q(
        \xmem_inst/mem[1][13] ), .QN(n1968) );
  DFF_X1 \xmem_inst/mem_reg[1][14]  ( .D(n838), .CK(clk), .Q(
        \xmem_inst/mem[1][14] ), .QN(n1969) );
  DFF_X1 \xmem_inst/mem_reg[1][15]  ( .D(n837), .CK(clk), .Q(
        \xmem_inst/mem[1][15] ), .QN(n1970) );
  DFF_X1 \xmem_inst/mem_reg[2][0]  ( .D(n836), .CK(clk), .Q(
        \xmem_inst/mem[2][0] ), .QN(n2052) );
  DFF_X1 \xmem_inst/mem_reg[2][1]  ( .D(n835), .CK(clk), .Q(
        \xmem_inst/mem[2][1] ), .QN(n2053) );
  DFF_X1 \xmem_inst/mem_reg[2][2]  ( .D(n834), .CK(clk), .Q(
        \xmem_inst/mem[2][2] ), .QN(n2054) );
  DFF_X1 \xmem_inst/mem_reg[2][3]  ( .D(n833), .CK(clk), .Q(
        \xmem_inst/mem[2][3] ), .QN(n2055) );
  DFF_X1 \xmem_inst/mem_reg[2][4]  ( .D(n832), .CK(clk), .Q(
        \xmem_inst/mem[2][4] ), .QN(n2056) );
  DFF_X1 \xmem_inst/mem_reg[2][5]  ( .D(n831), .CK(clk), .Q(
        \xmem_inst/mem[2][5] ), .QN(n2057) );
  DFF_X1 \xmem_inst/mem_reg[2][6]  ( .D(n830), .CK(clk), .Q(
        \xmem_inst/mem[2][6] ), .QN(n2058) );
  DFF_X1 \xmem_inst/mem_reg[2][7]  ( .D(n829), .CK(clk), .Q(
        \xmem_inst/mem[2][7] ), .QN(n2059) );
  DFF_X1 \xmem_inst/mem_reg[2][8]  ( .D(n828), .CK(clk), .Q(
        \xmem_inst/mem[2][8] ), .QN(n2060) );
  DFF_X1 \xmem_inst/mem_reg[2][9]  ( .D(n827), .CK(clk), .Q(
        \xmem_inst/mem[2][9] ), .QN(n2061) );
  DFF_X1 \xmem_inst/mem_reg[2][10]  ( .D(n826), .CK(clk), .Q(
        \xmem_inst/mem[2][10] ), .QN(n2062) );
  DFF_X1 \xmem_inst/mem_reg[2][11]  ( .D(n825), .CK(clk), .Q(
        \xmem_inst/mem[2][11] ), .QN(n2063) );
  DFF_X1 \xmem_inst/mem_reg[2][12]  ( .D(n824), .CK(clk), .Q(
        \xmem_inst/mem[2][12] ), .QN(n2064) );
  DFF_X1 \xmem_inst/mem_reg[2][13]  ( .D(n823), .CK(clk), .Q(
        \xmem_inst/mem[2][13] ), .QN(n2065) );
  DFF_X1 \xmem_inst/mem_reg[2][14]  ( .D(n822), .CK(clk), .Q(
        \xmem_inst/mem[2][14] ), .QN(n2066) );
  DFF_X1 \xmem_inst/mem_reg[2][15]  ( .D(n821), .CK(clk), .Q(
        \xmem_inst/mem[2][15] ), .QN(n2067) );
  DFF_X1 \xmem_inst/mem_reg[3][0]  ( .D(n820), .CK(clk), .Q(
        \xmem_inst/mem[3][0] ), .QN(n1971) );
  DFF_X1 \xmem_inst/mem_reg[3][1]  ( .D(n819), .CK(clk), .Q(
        \xmem_inst/mem[3][1] ), .QN(n1972) );
  DFF_X1 \xmem_inst/mem_reg[3][2]  ( .D(n818), .CK(clk), .Q(
        \xmem_inst/mem[3][2] ), .QN(n1973) );
  DFF_X1 \xmem_inst/mem_reg[3][3]  ( .D(n817), .CK(clk), .Q(
        \xmem_inst/mem[3][3] ), .QN(n1974) );
  DFF_X1 \xmem_inst/mem_reg[3][4]  ( .D(n816), .CK(clk), .Q(
        \xmem_inst/mem[3][4] ), .QN(n1975) );
  DFF_X1 \xmem_inst/mem_reg[3][5]  ( .D(n815), .CK(clk), .Q(
        \xmem_inst/mem[3][5] ), .QN(n1976) );
  DFF_X1 \xmem_inst/mem_reg[3][6]  ( .D(n814), .CK(clk), .Q(
        \xmem_inst/mem[3][6] ), .QN(n1977) );
  DFF_X1 \xmem_inst/mem_reg[3][7]  ( .D(n813), .CK(clk), .Q(
        \xmem_inst/mem[3][7] ), .QN(n1978) );
  DFF_X1 \xmem_inst/mem_reg[3][8]  ( .D(n812), .CK(clk), .Q(
        \xmem_inst/mem[3][8] ), .QN(n1979) );
  DFF_X1 \xmem_inst/mem_reg[3][9]  ( .D(n811), .CK(clk), .Q(
        \xmem_inst/mem[3][9] ), .QN(n1980) );
  DFF_X1 \xmem_inst/mem_reg[3][10]  ( .D(n810), .CK(clk), .Q(
        \xmem_inst/mem[3][10] ), .QN(n1981) );
  DFF_X1 \xmem_inst/mem_reg[3][11]  ( .D(n809), .CK(clk), .Q(
        \xmem_inst/mem[3][11] ), .QN(n1982) );
  DFF_X1 \xmem_inst/mem_reg[3][12]  ( .D(n808), .CK(clk), .Q(
        \xmem_inst/mem[3][12] ), .QN(n1983) );
  DFF_X1 \xmem_inst/mem_reg[3][13]  ( .D(n807), .CK(clk), .Q(
        \xmem_inst/mem[3][13] ), .QN(n1984) );
  DFF_X1 \xmem_inst/mem_reg[3][14]  ( .D(n806), .CK(clk), .Q(
        \xmem_inst/mem[3][14] ), .QN(n1985) );
  DFF_X1 \xmem_inst/mem_reg[3][15]  ( .D(n805), .CK(clk), .Q(
        \xmem_inst/mem[3][15] ), .QN(n1986) );
  DFF_X1 \xmem_inst/mem_reg[8][0]  ( .D(n740), .CK(clk), .Q(
        \xmem_inst/mem[8][0] ), .QN(n1875) );
  DFF_X1 \xmem_inst/mem_reg[8][1]  ( .D(n739), .CK(clk), .Q(
        \xmem_inst/mem[8][1] ), .QN(n1876) );
  DFF_X1 \xmem_inst/mem_reg[8][2]  ( .D(n738), .CK(clk), .Q(
        \xmem_inst/mem[8][2] ), .QN(n1877) );
  DFF_X1 \xmem_inst/mem_reg[8][3]  ( .D(n737), .CK(clk), .Q(
        \xmem_inst/mem[8][3] ), .QN(n1878) );
  DFF_X1 \xmem_inst/mem_reg[8][4]  ( .D(n736), .CK(clk), .Q(
        \xmem_inst/mem[8][4] ), .QN(n1879) );
  DFF_X1 \xmem_inst/mem_reg[8][5]  ( .D(n735), .CK(clk), .Q(
        \xmem_inst/mem[8][5] ), .QN(n1880) );
  DFF_X1 \xmem_inst/mem_reg[8][6]  ( .D(n734), .CK(clk), .Q(
        \xmem_inst/mem[8][6] ), .QN(n1881) );
  DFF_X1 \xmem_inst/mem_reg[8][7]  ( .D(n733), .CK(clk), .Q(
        \xmem_inst/mem[8][7] ), .QN(n1882) );
  DFF_X1 \xmem_inst/mem_reg[8][8]  ( .D(n732), .CK(clk), .Q(
        \xmem_inst/mem[8][8] ), .QN(n1883) );
  DFF_X1 \xmem_inst/mem_reg[8][9]  ( .D(n731), .CK(clk), .Q(
        \xmem_inst/mem[8][9] ), .QN(n1884) );
  DFF_X1 \xmem_inst/mem_reg[8][10]  ( .D(n730), .CK(clk), .Q(
        \xmem_inst/mem[8][10] ), .QN(n1885) );
  DFF_X1 \xmem_inst/mem_reg[8][11]  ( .D(n729), .CK(clk), .Q(
        \xmem_inst/mem[8][11] ), .QN(n1886) );
  DFF_X1 \xmem_inst/mem_reg[8][12]  ( .D(n728), .CK(clk), .Q(
        \xmem_inst/mem[8][12] ), .QN(n1887) );
  DFF_X1 \xmem_inst/mem_reg[8][13]  ( .D(n727), .CK(clk), .Q(
        \xmem_inst/mem[8][13] ), .QN(n1888) );
  DFF_X1 \xmem_inst/mem_reg[8][14]  ( .D(n726), .CK(clk), .Q(
        \xmem_inst/mem[8][14] ), .QN(n1889) );
  DFF_X1 \xmem_inst/mem_reg[8][15]  ( .D(n725), .CK(clk), .Q(
        \xmem_inst/mem[8][15] ), .QN(n1890) );
  DFF_X1 \xmem_inst/mem_reg[9][0]  ( .D(n724), .CK(clk), .Q(
        \xmem_inst/mem[9][0] ), .QN(n1891) );
  DFF_X1 \xmem_inst/mem_reg[9][1]  ( .D(n723), .CK(clk), .Q(
        \xmem_inst/mem[9][1] ), .QN(n1892) );
  DFF_X1 \xmem_inst/mem_reg[9][2]  ( .D(n722), .CK(clk), .Q(
        \xmem_inst/mem[9][2] ), .QN(n1893) );
  DFF_X1 \xmem_inst/mem_reg[9][3]  ( .D(n721), .CK(clk), .Q(
        \xmem_inst/mem[9][3] ), .QN(n1894) );
  DFF_X1 \xmem_inst/mem_reg[9][4]  ( .D(n720), .CK(clk), .Q(
        \xmem_inst/mem[9][4] ), .QN(n1895) );
  DFF_X1 \xmem_inst/mem_reg[9][5]  ( .D(n719), .CK(clk), .Q(
        \xmem_inst/mem[9][5] ), .QN(n1896) );
  DFF_X1 \xmem_inst/mem_reg[9][6]  ( .D(n718), .CK(clk), .Q(
        \xmem_inst/mem[9][6] ), .QN(n1897) );
  DFF_X1 \xmem_inst/mem_reg[9][7]  ( .D(n717), .CK(clk), .Q(
        \xmem_inst/mem[9][7] ), .QN(n1898) );
  DFF_X1 \xmem_inst/mem_reg[9][8]  ( .D(n716), .CK(clk), .Q(
        \xmem_inst/mem[9][8] ), .QN(n1899) );
  DFF_X1 \xmem_inst/mem_reg[9][9]  ( .D(n715), .CK(clk), .Q(
        \xmem_inst/mem[9][9] ), .QN(n1900) );
  DFF_X1 \xmem_inst/mem_reg[9][10]  ( .D(n714), .CK(clk), .Q(
        \xmem_inst/mem[9][10] ), .QN(n1901) );
  DFF_X1 \xmem_inst/mem_reg[9][11]  ( .D(n713), .CK(clk), .Q(
        \xmem_inst/mem[9][11] ), .QN(n1902) );
  DFF_X1 \xmem_inst/mem_reg[9][12]  ( .D(n712), .CK(clk), .Q(
        \xmem_inst/mem[9][12] ), .QN(n1903) );
  DFF_X1 \xmem_inst/mem_reg[9][13]  ( .D(n711), .CK(clk), .Q(
        \xmem_inst/mem[9][13] ), .QN(n1904) );
  DFF_X1 \xmem_inst/mem_reg[9][14]  ( .D(n710), .CK(clk), .Q(
        \xmem_inst/mem[9][14] ), .QN(n1905) );
  DFF_X1 \xmem_inst/mem_reg[9][15]  ( .D(n709), .CK(clk), .Q(
        \xmem_inst/mem[9][15] ), .QN(n1906) );
  DFF_X1 \xmem_inst/mem_reg[10][0]  ( .D(n708), .CK(clk), .Q(
        \xmem_inst/mem[10][0] ), .QN(n1907) );
  DFF_X1 \xmem_inst/mem_reg[10][1]  ( .D(n707), .CK(clk), .Q(
        \xmem_inst/mem[10][1] ), .QN(n1908) );
  DFF_X1 \xmem_inst/mem_reg[10][2]  ( .D(n706), .CK(clk), .Q(
        \xmem_inst/mem[10][2] ), .QN(n1909) );
  DFF_X1 \xmem_inst/mem_reg[10][3]  ( .D(n705), .CK(clk), .Q(
        \xmem_inst/mem[10][3] ), .QN(n1910) );
  DFF_X1 \xmem_inst/mem_reg[10][4]  ( .D(n704), .CK(clk), .Q(
        \xmem_inst/mem[10][4] ), .QN(n1911) );
  DFF_X1 \xmem_inst/mem_reg[10][5]  ( .D(n703), .CK(clk), .Q(
        \xmem_inst/mem[10][5] ), .QN(n1912) );
  DFF_X1 \xmem_inst/mem_reg[10][6]  ( .D(n702), .CK(clk), .Q(
        \xmem_inst/mem[10][6] ), .QN(n1913) );
  DFF_X1 \xmem_inst/mem_reg[10][7]  ( .D(n701), .CK(clk), .Q(
        \xmem_inst/mem[10][7] ), .QN(n1914) );
  DFF_X1 \xmem_inst/mem_reg[10][8]  ( .D(n700), .CK(clk), .Q(
        \xmem_inst/mem[10][8] ), .QN(n1915) );
  DFF_X1 \xmem_inst/mem_reg[10][9]  ( .D(n699), .CK(clk), .Q(
        \xmem_inst/mem[10][9] ), .QN(n1916) );
  DFF_X1 \xmem_inst/mem_reg[10][10]  ( .D(n698), .CK(clk), .Q(
        \xmem_inst/mem[10][10] ), .QN(n1917) );
  DFF_X1 \xmem_inst/mem_reg[10][11]  ( .D(n697), .CK(clk), .Q(
        \xmem_inst/mem[10][11] ), .QN(n1918) );
  DFF_X1 \xmem_inst/mem_reg[10][12]  ( .D(n696), .CK(clk), .Q(
        \xmem_inst/mem[10][12] ), .QN(n1919) );
  DFF_X1 \xmem_inst/mem_reg[10][13]  ( .D(n695), .CK(clk), .Q(
        \xmem_inst/mem[10][13] ), .QN(n1920) );
  DFF_X1 \xmem_inst/mem_reg[10][14]  ( .D(n694), .CK(clk), .Q(
        \xmem_inst/mem[10][14] ), .QN(n1921) );
  DFF_X1 \xmem_inst/mem_reg[10][15]  ( .D(n693), .CK(clk), .Q(
        \xmem_inst/mem[10][15] ), .QN(n1922) );
  DFF_X1 \xmem_inst/mem_reg[11][0]  ( .D(n692), .CK(clk), .Q(
        \xmem_inst/mem[11][0] ), .QN(n1923) );
  DFF_X1 \xmem_inst/mem_reg[11][1]  ( .D(n691), .CK(clk), .Q(
        \xmem_inst/mem[11][1] ), .QN(n1924) );
  DFF_X1 \xmem_inst/mem_reg[11][2]  ( .D(n690), .CK(clk), .Q(
        \xmem_inst/mem[11][2] ), .QN(n1925) );
  DFF_X1 \xmem_inst/mem_reg[11][3]  ( .D(n689), .CK(clk), .Q(
        \xmem_inst/mem[11][3] ), .QN(n1926) );
  DFF_X1 \xmem_inst/mem_reg[11][4]  ( .D(n688), .CK(clk), .Q(
        \xmem_inst/mem[11][4] ), .QN(n1927) );
  DFF_X1 \xmem_inst/mem_reg[11][5]  ( .D(n687), .CK(clk), .Q(
        \xmem_inst/mem[11][5] ), .QN(n1928) );
  DFF_X1 \xmem_inst/mem_reg[11][6]  ( .D(n686), .CK(clk), .Q(
        \xmem_inst/mem[11][6] ), .QN(n1929) );
  DFF_X1 \xmem_inst/mem_reg[11][7]  ( .D(n685), .CK(clk), .Q(
        \xmem_inst/mem[11][7] ), .QN(n1930) );
  DFF_X1 \xmem_inst/mem_reg[11][8]  ( .D(n684), .CK(clk), .Q(
        \xmem_inst/mem[11][8] ), .QN(n1931) );
  DFF_X1 \xmem_inst/mem_reg[11][9]  ( .D(n683), .CK(clk), .Q(
        \xmem_inst/mem[11][9] ), .QN(n1932) );
  DFF_X1 \xmem_inst/mem_reg[11][10]  ( .D(n682), .CK(clk), .Q(
        \xmem_inst/mem[11][10] ), .QN(n1933) );
  DFF_X1 \xmem_inst/mem_reg[11][11]  ( .D(n681), .CK(clk), .Q(
        \xmem_inst/mem[11][11] ), .QN(n1934) );
  DFF_X1 \xmem_inst/mem_reg[11][12]  ( .D(n680), .CK(clk), .Q(
        \xmem_inst/mem[11][12] ), .QN(n1935) );
  DFF_X1 \xmem_inst/mem_reg[11][13]  ( .D(n679), .CK(clk), .Q(
        \xmem_inst/mem[11][13] ), .QN(n1936) );
  DFF_X1 \xmem_inst/mem_reg[11][14]  ( .D(n678), .CK(clk), .Q(
        \xmem_inst/mem[11][14] ), .QN(n1937) );
  DFF_X1 \xmem_inst/mem_reg[11][15]  ( .D(n677), .CK(clk), .Q(
        \xmem_inst/mem[11][15] ), .QN(n1938) );
  DFF_X1 \xmem_inst/mem_reg[15][0]  ( .D(n628), .CK(clk), .Q(
        \xmem_inst/mem[15][0] ), .QN(n2019) );
  DFF_X1 \xmem_inst/mem_reg[15][1]  ( .D(n627), .CK(clk), .Q(
        \xmem_inst/mem[15][1] ), .QN(n2020) );
  DFF_X1 \xmem_inst/mem_reg[15][2]  ( .D(n626), .CK(clk), .Q(
        \xmem_inst/mem[15][2] ), .QN(n2021) );
  DFF_X1 \xmem_inst/mem_reg[15][3]  ( .D(n625), .CK(clk), .Q(
        \xmem_inst/mem[15][3] ), .QN(n2022) );
  DFF_X1 \xmem_inst/mem_reg[15][4]  ( .D(n624), .CK(clk), .Q(
        \xmem_inst/mem[15][4] ), .QN(n2023) );
  DFF_X1 \xmem_inst/mem_reg[15][5]  ( .D(n623), .CK(clk), .Q(
        \xmem_inst/mem[15][5] ), .QN(n2024) );
  DFF_X1 \xmem_inst/mem_reg[15][6]  ( .D(n622), .CK(clk), .Q(
        \xmem_inst/mem[15][6] ), .QN(n2025) );
  DFF_X1 \xmem_inst/mem_reg[15][7]  ( .D(n621), .CK(clk), .Q(
        \xmem_inst/mem[15][7] ), .QN(n2026) );
  DFF_X1 \xmem_inst/mem_reg[15][8]  ( .D(n620), .CK(clk), .Q(
        \xmem_inst/mem[15][8] ), .QN(n2027) );
  DFF_X1 \xmem_inst/mem_reg[15][9]  ( .D(n619), .CK(clk), .Q(
        \xmem_inst/mem[15][9] ), .QN(n2028) );
  DFF_X1 \xmem_inst/mem_reg[15][10]  ( .D(n618), .CK(clk), .Q(
        \xmem_inst/mem[15][10] ), .QN(n2029) );
  DFF_X1 \xmem_inst/mem_reg[15][11]  ( .D(n617), .CK(clk), .Q(
        \xmem_inst/mem[15][11] ), .QN(n2030) );
  DFF_X1 \xmem_inst/mem_reg[15][12]  ( .D(n616), .CK(clk), .Q(
        \xmem_inst/mem[15][12] ), .QN(n2031) );
  DFF_X1 \xmem_inst/mem_reg[15][13]  ( .D(n615), .CK(clk), .Q(
        \xmem_inst/mem[15][13] ), .QN(n2032) );
  DFF_X1 \xmem_inst/mem_reg[15][14]  ( .D(n614), .CK(clk), .Q(
        \xmem_inst/mem[15][14] ), .QN(n2033) );
  DFF_X1 \xmem_inst/mem_reg[15][15]  ( .D(n613), .CK(clk), .Q(
        \xmem_inst/mem[15][15] ), .QN(n2034) );
  DFF_X1 \ctrl_conv_output_inst/conv_start_accum_reg  ( .D(n2133), .CK(clk), 
        .Q(\ctrl_conv_output_inst/conv_start_accum ) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[0]  ( .D(n595), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [0]), .QN(n1868) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[1]  ( .D(n594), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [1]), .QN(n1865) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[2]  ( .D(n593), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [2]), .QN(n1866) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[3]  ( .D(n592), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [3]), .QN(n1864) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[4]  ( .D(n591), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [4]), .QN(n1869) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[5]  ( .D(n590), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [5]), .QN(n1871) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[6]  ( .D(n589), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [6]), .QN(n1867) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[7]  ( .D(n588), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [7]), .QN(n1872) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[8]  ( .D(n587), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [8]), .QN(n1843) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[9]  ( .D(n586), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [9]), .QN(n1844) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[10]  ( .D(n585), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [10]), .QN(n1845) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[11]  ( .D(n584), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [11]), .QN(n1873) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[12]  ( .D(n583), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [12]), .QN(n1846) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[13]  ( .D(n582), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [13]), .QN(n1874) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[14]  ( .D(n581), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [14]), .QN(n1847) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[2]  ( .D(n609), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [2]), .QN(n2120) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[4]  ( .D(n607), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [4]), .QN(n2122) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[5]  ( .D(n606), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [5]), .QN(n2123) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[10]  ( .D(n601), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [10]), .QN(n2128) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[11]  ( .D(n600), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [11]), .QN(n2129) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[13]  ( .D(n598), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [13]), .QN(n2131) );
  DFF_X1 \fmem_addr_reg[0]  ( .D(n578), .CK(clk), .Q(\fmem_inst/N14 ), .QN(
        n1834) );
  DFF_X1 \fmem_inst/z_reg[0]  ( .D(\fmem_inst/N12 ), .CK(clk), .Q(n1816), .QN(
        n1823) );
  DFF_X1 \xmem_inst/data_out_reg[11]  ( .D(\xmem_inst/N18 ), .CK(clk), .Q(
        xmem_data[11]), .QN(n1827) );
  DFF_X1 \xmem_inst/data_out_reg[0]  ( .D(\xmem_inst/N29 ), .CK(clk), .Q(
        xmem_data[0]), .QN(n1824) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[3]  ( .D(n878), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [3]) );
  DFF_X1 \fmem_addr_reg[1]  ( .D(n579), .CK(clk), .Q(\fmem_inst/N12 ) );
  DFF_X1 \xmem_inst/data_out_reg[1]  ( .D(\xmem_inst/N28 ), .CK(clk), .QN(
        n1830) );
  DFF_X1 \xmem_inst/data_out_reg[4]  ( .D(\xmem_inst/N25 ), .CK(clk), .QN(
        n1829) );
  DFF_X1 \xmem_inst/data_out_reg[5]  ( .D(\xmem_inst/N24 ), .CK(clk), .QN(
        n1825) );
  DFF_X1 \xmem_inst/data_out_reg[15]  ( .D(\xmem_inst/N14 ), .CK(clk), .QN(
        n1826) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[15]  ( .D(n596), .CK(clk), .QN(n1822)
         );
  DFF_X1 \mac_unit_inst/adder_reg_reg[15]  ( .D(n580), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [15]), .QN(n1839) );
  DFF_X2 \mac_unit_inst/x_mult_f_reg_reg[14]  ( .D(n597), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [14]), .QN(n2132) );
  DFF_X1 \fmem_inst/z_reg[6]  ( .D(\fmem_inst/N13 ), .CK(clk), .Q(n1821), .QN(
        n1828) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[12]  ( .D(n599), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [12]), .QN(n2130) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[0]  ( .D(n611), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [0]), .QN(n2118) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[9]  ( .D(n602), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [9]), .QN(n2127) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[8]  ( .D(n603), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [8]), .QN(n2126) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[6]  ( .D(n605), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [6]), .QN(n2124) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[7]  ( .D(n604), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [7]), .QN(n2125) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[3]  ( .D(n608), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [3]), .QN(n2121) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[1]  ( .D(n610), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [1]), .QN(n2119) );
  BUF_X1 U919 ( .A(n1823), .Z(n1283) );
  AND2_X1 U920 ( .A1(n1821), .A2(xmem_data[14]), .ZN(n1250) );
  NOR2_X1 U921 ( .A1(n882), .A2(n1832), .ZN(n1374) );
  AND2_X1 U922 ( .A1(n1345), .A2(n1344), .ZN(n1634) );
  OR2_X1 U923 ( .A1(n1345), .A2(n1344), .ZN(n1636) );
  NOR2_X1 U924 ( .A1(n903), .A2(n1411), .ZN(n880) );
  NAND2_X1 U925 ( .A1(n1477), .A2(n1476), .ZN(n1589) );
  OR2_X1 U926 ( .A1(n1255), .A2(n1254), .ZN(n1598) );
  INV_X1 U927 ( .A(n1770), .ZN(n1769) );
  INV_X1 U928 ( .A(n1780), .ZN(n1781) );
  INV_X1 U929 ( .A(n1757), .ZN(n1758) );
  INV_X1 U930 ( .A(n1808), .ZN(n1810) );
  INV_X1 U931 ( .A(n1766), .ZN(n1765) );
  NAND2_X1 U932 ( .A1(n1786), .A2(n1735), .ZN(n1808) );
  NAND2_X1 U933 ( .A1(n1786), .A2(n1779), .ZN(n1780) );
  INV_X1 U934 ( .A(n1755), .ZN(n1754) );
  INV_X1 U935 ( .A(n1792), .ZN(n1791) );
  INV_X1 U936 ( .A(n1784), .ZN(n1783) );
  INV_X1 U937 ( .A(n1787), .ZN(n1788) );
  INV_X1 U938 ( .A(n1774), .ZN(n1775) );
  INV_X1 U939 ( .A(n1772), .ZN(n1771) );
  INV_X1 U940 ( .A(n1760), .ZN(n1759) );
  INV_X1 U941 ( .A(n1748), .ZN(n1747) );
  INV_X1 U942 ( .A(n1750), .ZN(n1751) );
  INV_X1 U943 ( .A(n1762), .ZN(n1763) );
  NAND2_X1 U944 ( .A1(n1786), .A2(n1756), .ZN(n1757) );
  INV_X1 U945 ( .A(n1778), .ZN(n1777) );
  NAND2_X1 U946 ( .A1(n1786), .A2(n1761), .ZN(n1762) );
  NAND2_X1 U947 ( .A1(n1786), .A2(n1773), .ZN(n1774) );
  NAND2_X1 U948 ( .A1(n1786), .A2(n1785), .ZN(n1787) );
  NAND2_X1 U949 ( .A1(n1786), .A2(n1749), .ZN(n1750) );
  OR2_X1 U950 ( .A1(n1123), .A2(n1764), .ZN(n1767) );
  OR2_X1 U951 ( .A1(n1283), .A2(n1826), .ZN(n1201) );
  AND2_X1 U952 ( .A1(n1821), .A2(xmem_data[12]), .ZN(n1271) );
  BUF_X2 U953 ( .A(n1828), .Z(n881) );
  BUF_X2 U954 ( .A(n1828), .Z(n882) );
  INV_X1 U955 ( .A(n1310), .ZN(n1294) );
  NAND2_X1 U956 ( .A1(n1333), .A2(n1310), .ZN(n1318) );
  NAND2_X1 U957 ( .A1(n1238), .A2(n1237), .ZN(n1441) );
  NAND2_X1 U958 ( .A1(n1246), .A2(n1244), .ZN(n1237) );
  OR2_X1 U959 ( .A1(n1320), .A2(n1323), .ZN(n1321) );
  XNOR2_X1 U960 ( .A(n1301), .B(n1300), .ZN(n1322) );
  AND2_X1 U961 ( .A1(n1336), .A2(n1374), .ZN(n1344) );
  CLKBUF_X1 U962 ( .A(n1637), .Z(n885) );
  CLKBUF_X1 U963 ( .A(n1642), .Z(n893) );
  OR2_X1 U964 ( .A1(n1349), .A2(n1348), .ZN(n1649) );
  INV_X1 U965 ( .A(n1634), .ZN(n1635) );
  OR2_X1 U966 ( .A1(n1326), .A2(n1826), .ZN(n1234) );
  NAND2_X1 U967 ( .A1(n1177), .A2(n1176), .ZN(n1178) );
  INV_X1 U968 ( .A(n1373), .ZN(n1303) );
  NAND2_X1 U969 ( .A1(n1364), .A2(n1363), .ZN(n1365) );
  NAND2_X1 U970 ( .A1(n1362), .A2(n1361), .ZN(n1363) );
  OR2_X1 U971 ( .A1(n1362), .A2(n1361), .ZN(n1359) );
  XOR2_X1 U972 ( .A(n1444), .B(n1443), .Z(n1242) );
  NAND2_X1 U973 ( .A1(n1301), .A2(n1284), .ZN(n1286) );
  NAND2_X1 U974 ( .A1(n1314), .A2(n1313), .ZN(n1391) );
  NAND2_X1 U975 ( .A1(n1382), .A2(n1380), .ZN(n1313) );
  OAI21_X1 U976 ( .B1(n1382), .B2(n1380), .A(n896), .ZN(n1314) );
  CLKBUF_X1 U977 ( .A(n1381), .Z(n896) );
  NAND2_X1 U978 ( .A1(n1306), .A2(n1305), .ZN(n1382) );
  NAND2_X1 U979 ( .A1(n1374), .A2(n1373), .ZN(n1305) );
  NAND2_X1 U980 ( .A1(n1376), .A2(n1304), .ZN(n1306) );
  NAND2_X1 U981 ( .A1(n1337), .A2(n1303), .ZN(n1304) );
  NAND2_X1 U982 ( .A1(n1320), .A2(n1323), .ZN(n1324) );
  NAND2_X1 U983 ( .A1(n1322), .A2(n1321), .ZN(n1325) );
  XNOR2_X1 U984 ( .A(n1328), .B(n1361), .ZN(n1329) );
  XNOR2_X1 U985 ( .A(n1222), .B(n1221), .ZN(n1224) );
  CLKBUF_X1 U986 ( .A(n1697), .Z(n900) );
  NAND2_X1 U987 ( .A1(s_ready_x), .A2(s_valid_x), .ZN(n1768) );
  OR2_X1 U988 ( .A1(n1768), .A2(n1752), .ZN(n1789) );
  INV_X1 U989 ( .A(n1768), .ZN(n1786) );
  OR2_X1 U990 ( .A1(n1768), .A2(n1746), .ZN(n1782) );
  CLKBUF_X1 U991 ( .A(n1651), .Z(n1652) );
  CLKBUF_X1 U992 ( .A(n1670), .Z(n883) );
  AND2_X1 U993 ( .A1(n1167), .A2(n1165), .ZN(n1477) );
  CLKBUF_X1 U994 ( .A(n1593), .Z(n892) );
  INV_X1 U995 ( .A(n1127), .ZN(n1123) );
  CLKBUF_X1 U996 ( .A(n1656), .Z(n1661) );
  NAND2_X1 U997 ( .A1(n1636), .A2(n1635), .ZN(n1638) );
  AND2_X1 U998 ( .A1(n1821), .A2(xmem_data[10]), .ZN(n1298) );
  AND2_X1 U999 ( .A1(n1821), .A2(xmem_data[6]), .ZN(n1354) );
  XNOR2_X1 U1000 ( .A(n1224), .B(n1223), .ZN(n1417) );
  AND2_X1 U1001 ( .A1(n1338), .A2(xmem_data[0]), .ZN(n884) );
  NAND2_X1 U1002 ( .A1(n1355), .A2(n1274), .ZN(n1188) );
  OR2_X1 U1003 ( .A1(n1274), .A2(n1355), .ZN(n1187) );
  AND2_X1 U1004 ( .A1(n1821), .A2(xmem_data[11]), .ZN(n886) );
  XOR2_X1 U1005 ( .A(n1281), .B(n1282), .Z(n887) );
  XOR2_X1 U1006 ( .A(n1280), .B(n887), .Z(n1316) );
  NAND2_X1 U1007 ( .A1(n1280), .A2(n1281), .ZN(n888) );
  NAND2_X1 U1008 ( .A1(n1280), .A2(n1282), .ZN(n889) );
  NAND2_X1 U1009 ( .A1(n1281), .A2(n1282), .ZN(n890) );
  NAND3_X1 U1010 ( .A1(n888), .A2(n889), .A3(n890), .ZN(n1276) );
  NOR2_X1 U1011 ( .A1(n1427), .A2(n1426), .ZN(n891) );
  AND2_X1 U1012 ( .A1(n1821), .A2(xmem_data[11]), .ZN(n1280) );
  AOI21_X1 U1013 ( .B1(n1636), .B2(n1637), .A(n1634), .ZN(n894) );
  AND2_X1 U1014 ( .A1(n1816), .A2(xmem_data[12]), .ZN(n1282) );
  BUF_X1 U1015 ( .A(n1231), .Z(n895) );
  NAND2_X1 U1016 ( .A1(n1180), .A2(n1179), .ZN(n897) );
  NOR2_X1 U1017 ( .A1(n1394), .A2(n1393), .ZN(n898) );
  NOR2_X1 U1018 ( .A1(n1394), .A2(n1393), .ZN(n1689) );
  NOR2_X1 U1019 ( .A1(n1398), .A2(n1397), .ZN(n899) );
  NAND2_X1 U1020 ( .A1(n1360), .A2(n1359), .ZN(n1364) );
  XNOR2_X1 U1021 ( .A(n1360), .B(n1329), .ZN(n1349) );
  INV_X1 U1022 ( .A(n1707), .ZN(n901) );
  NAND2_X1 U1023 ( .A1(n1604), .A2(n1603), .ZN(n902) );
  FA_X1 U1024 ( .A(n897), .B(n1219), .CI(n1218), .CO(n903) );
  BUF_X1 U1025 ( .A(n1620), .Z(n904) );
  BUF_X1 U1026 ( .A(n1620), .Z(n905) );
  AND2_X1 U1027 ( .A1(n1415), .A2(n1414), .ZN(n910) );
  XOR2_X1 U1028 ( .A(n1451), .B(n1450), .Z(n912) );
  XOR2_X1 U1029 ( .A(n1434), .B(n1433), .Z(n913) );
  XOR2_X1 U1030 ( .A(n1440), .B(n1439), .Z(n914) );
  NOR2_X1 U1031 ( .A1(n1444), .A2(n1443), .ZN(n915) );
  NOR2_X1 U1032 ( .A1(n1434), .A2(n1433), .ZN(n916) );
  OR2_X1 U1033 ( .A1(n1439), .A2(n1440), .ZN(n917) );
  NAND2_X1 U1034 ( .A1(n1833), .A2(n1838), .ZN(n1746) );
  NAND2_X1 U1035 ( .A1(xmem_addr[2]), .A2(xmem_addr[3]), .ZN(n1790) );
  NOR2_X2 U1036 ( .A1(n1746), .A2(n1790), .ZN(n1098) );
  NAND2_X1 U1037 ( .A1(xmem_addr[0]), .A2(n1838), .ZN(n1741) );
  NOR2_X2 U1038 ( .A1(n1741), .A2(n1790), .ZN(n1785) );
  AOI22_X1 U1039 ( .A1(n1098), .A2(\xmem_inst/mem[12][3] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][3] ), .ZN(n921) );
  NAND2_X1 U1040 ( .A1(xmem_addr[1]), .A2(n1833), .ZN(n1752) );
  NOR2_X2 U1041 ( .A1(n1752), .A2(n1790), .ZN(n1099) );
  NOR2_X1 U1042 ( .A1(n1833), .A2(n1838), .ZN(n1127) );
  NOR2_X2 U1043 ( .A1(n1123), .A2(n1790), .ZN(n1735) );
  AOI22_X1 U1044 ( .A1(n1099), .A2(\xmem_inst/mem[14][3] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][3] ), .ZN(n920) );
  NAND2_X1 U1045 ( .A1(n1835), .A2(n1842), .ZN(n1753) );
  NOR2_X2 U1046 ( .A1(n1746), .A2(n1753), .ZN(n1100) );
  NOR2_X2 U1047 ( .A1(n1741), .A2(n1753), .ZN(n1749) );
  AOI22_X1 U1048 ( .A1(n1100), .A2(\xmem_inst/mem[0][3] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][3] ), .ZN(n919) );
  NOR2_X2 U1049 ( .A1(n1752), .A2(n1753), .ZN(n1101) );
  NOR2_X2 U1050 ( .A1(n1123), .A2(n1753), .ZN(n1756) );
  AOI22_X1 U1051 ( .A1(n1101), .A2(\xmem_inst/mem[2][3] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][3] ), .ZN(n918) );
  NAND4_X1 U1052 ( .A1(n921), .A2(n920), .A3(n919), .A4(n918), .ZN(n929) );
  NAND2_X1 U1053 ( .A1(n1842), .A2(xmem_addr[2]), .ZN(n1764) );
  NOR2_X2 U1054 ( .A1(n1764), .A2(n1746), .ZN(n1106) );
  NOR2_X2 U1055 ( .A1(n1764), .A2(n1741), .ZN(n1761) );
  AOI22_X1 U1056 ( .A1(n1106), .A2(\xmem_inst/mem[4][3] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][3] ), .ZN(n922) );
  OAI21_X1 U1057 ( .B1(n1767), .B2(n1851), .A(n922), .ZN(n928) );
  NAND2_X1 U1058 ( .A1(xmem_addr[3]), .A2(n1835), .ZN(n1776) );
  NOR2_X2 U1059 ( .A1(n1123), .A2(n1776), .ZN(n1779) );
  NAND2_X1 U1060 ( .A1(n1779), .A2(\xmem_inst/mem[11][3] ), .ZN(n926) );
  NOR2_X2 U1061 ( .A1(n1764), .A2(n1752), .ZN(n1109) );
  NOR2_X2 U1062 ( .A1(n1776), .A2(n1746), .ZN(n1108) );
  AOI22_X1 U1063 ( .A1(n1109), .A2(\xmem_inst/mem[6][3] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][3] ), .ZN(n925) );
  NOR2_X2 U1064 ( .A1(n1776), .A2(n1741), .ZN(n1773) );
  NAND2_X1 U1065 ( .A1(n1773), .A2(\xmem_inst/mem[9][3] ), .ZN(n924) );
  NOR2_X2 U1066 ( .A1(n1776), .A2(n1752), .ZN(n1110) );
  NAND2_X1 U1067 ( .A1(n1110), .A2(\xmem_inst/mem[10][3] ), .ZN(n923) );
  NAND4_X1 U1068 ( .A1(n926), .A2(n925), .A3(n924), .A4(n923), .ZN(n927) );
  OR3_X1 U1069 ( .A1(n929), .A2(n928), .A3(n927), .ZN(\xmem_inst/N26 ) );
  AOI22_X1 U1070 ( .A1(n1098), .A2(\xmem_inst/mem[12][15] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][15] ), .ZN(n933) );
  AOI22_X1 U1071 ( .A1(n1099), .A2(\xmem_inst/mem[14][15] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][15] ), .ZN(n932) );
  AOI22_X1 U1072 ( .A1(n1100), .A2(\xmem_inst/mem[0][15] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][15] ), .ZN(n931) );
  AOI22_X1 U1073 ( .A1(n1101), .A2(\xmem_inst/mem[2][15] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][15] ), .ZN(n930) );
  NAND4_X1 U1074 ( .A1(n933), .A2(n932), .A3(n931), .A4(n930), .ZN(n941) );
  AOI22_X1 U1075 ( .A1(n1106), .A2(\xmem_inst/mem[4][15] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][15] ), .ZN(n934) );
  OAI21_X1 U1076 ( .B1(n1767), .B2(n1863), .A(n934), .ZN(n940) );
  NAND2_X1 U1077 ( .A1(n1779), .A2(\xmem_inst/mem[11][15] ), .ZN(n938) );
  AOI22_X1 U1078 ( .A1(n1109), .A2(\xmem_inst/mem[6][15] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][15] ), .ZN(n937) );
  NAND2_X1 U1079 ( .A1(n1773), .A2(\xmem_inst/mem[9][15] ), .ZN(n936) );
  NAND2_X1 U1080 ( .A1(n1110), .A2(\xmem_inst/mem[10][15] ), .ZN(n935) );
  NAND4_X1 U1081 ( .A1(n938), .A2(n937), .A3(n936), .A4(n935), .ZN(n939) );
  OR3_X1 U1082 ( .A1(n941), .A2(n940), .A3(n939), .ZN(\xmem_inst/N14 ) );
  AOI22_X1 U1083 ( .A1(n1098), .A2(\xmem_inst/mem[12][4] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][4] ), .ZN(n945) );
  AOI22_X1 U1084 ( .A1(n1099), .A2(\xmem_inst/mem[14][4] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][4] ), .ZN(n944) );
  AOI22_X1 U1085 ( .A1(n1100), .A2(\xmem_inst/mem[0][4] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][4] ), .ZN(n943) );
  AOI22_X1 U1086 ( .A1(n1101), .A2(\xmem_inst/mem[2][4] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][4] ), .ZN(n942) );
  NAND4_X1 U1087 ( .A1(n945), .A2(n944), .A3(n943), .A4(n942), .ZN(n953) );
  AOI22_X1 U1088 ( .A1(n1106), .A2(\xmem_inst/mem[4][4] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][4] ), .ZN(n946) );
  OAI21_X1 U1089 ( .B1(n1767), .B2(n1852), .A(n946), .ZN(n952) );
  NAND2_X1 U1090 ( .A1(n1779), .A2(\xmem_inst/mem[11][4] ), .ZN(n950) );
  AOI22_X1 U1091 ( .A1(n1109), .A2(\xmem_inst/mem[6][4] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][4] ), .ZN(n949) );
  NAND2_X1 U1092 ( .A1(n1773), .A2(\xmem_inst/mem[9][4] ), .ZN(n948) );
  NAND2_X1 U1093 ( .A1(n1110), .A2(\xmem_inst/mem[10][4] ), .ZN(n947) );
  NAND4_X1 U1094 ( .A1(n950), .A2(n949), .A3(n948), .A4(n947), .ZN(n951) );
  OR3_X1 U1095 ( .A1(n953), .A2(n952), .A3(n951), .ZN(\xmem_inst/N25 ) );
  AOI22_X1 U1096 ( .A1(n1098), .A2(\xmem_inst/mem[12][5] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][5] ), .ZN(n957) );
  AOI22_X1 U1097 ( .A1(n1099), .A2(\xmem_inst/mem[14][5] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][5] ), .ZN(n956) );
  AOI22_X1 U1098 ( .A1(n1100), .A2(\xmem_inst/mem[0][5] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][5] ), .ZN(n955) );
  AOI22_X1 U1099 ( .A1(n1101), .A2(\xmem_inst/mem[2][5] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][5] ), .ZN(n954) );
  NAND4_X1 U1100 ( .A1(n957), .A2(n956), .A3(n955), .A4(n954), .ZN(n965) );
  AOI22_X1 U1101 ( .A1(n1106), .A2(\xmem_inst/mem[4][5] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][5] ), .ZN(n958) );
  OAI21_X1 U1102 ( .B1(n1767), .B2(n1853), .A(n958), .ZN(n964) );
  NAND2_X1 U1103 ( .A1(n1779), .A2(\xmem_inst/mem[11][5] ), .ZN(n962) );
  AOI22_X1 U1104 ( .A1(n1109), .A2(\xmem_inst/mem[6][5] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][5] ), .ZN(n961) );
  NAND2_X1 U1105 ( .A1(n1773), .A2(\xmem_inst/mem[9][5] ), .ZN(n960) );
  NAND2_X1 U1106 ( .A1(n1110), .A2(\xmem_inst/mem[10][5] ), .ZN(n959) );
  NAND4_X1 U1107 ( .A1(n962), .A2(n961), .A3(n960), .A4(n959), .ZN(n963) );
  OR3_X1 U1108 ( .A1(n965), .A2(n964), .A3(n963), .ZN(\xmem_inst/N24 ) );
  AOI22_X1 U1109 ( .A1(n1098), .A2(\xmem_inst/mem[12][6] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][6] ), .ZN(n969) );
  AOI22_X1 U1110 ( .A1(n1099), .A2(\xmem_inst/mem[14][6] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][6] ), .ZN(n968) );
  AOI22_X1 U1111 ( .A1(n1100), .A2(\xmem_inst/mem[0][6] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][6] ), .ZN(n967) );
  AOI22_X1 U1112 ( .A1(n1101), .A2(\xmem_inst/mem[2][6] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][6] ), .ZN(n966) );
  NAND4_X1 U1113 ( .A1(n969), .A2(n968), .A3(n967), .A4(n966), .ZN(n977) );
  AOI22_X1 U1114 ( .A1(n1106), .A2(\xmem_inst/mem[4][6] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][6] ), .ZN(n970) );
  OAI21_X1 U1115 ( .B1(n1767), .B2(n1854), .A(n970), .ZN(n976) );
  NAND2_X1 U1116 ( .A1(n1779), .A2(\xmem_inst/mem[11][6] ), .ZN(n974) );
  AOI22_X1 U1117 ( .A1(n1109), .A2(\xmem_inst/mem[6][6] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][6] ), .ZN(n973) );
  NAND2_X1 U1118 ( .A1(n1773), .A2(\xmem_inst/mem[9][6] ), .ZN(n972) );
  NAND2_X1 U1119 ( .A1(n1110), .A2(\xmem_inst/mem[10][6] ), .ZN(n971) );
  NAND4_X1 U1120 ( .A1(n974), .A2(n973), .A3(n972), .A4(n971), .ZN(n975) );
  OR3_X1 U1121 ( .A1(n977), .A2(n976), .A3(n975), .ZN(\xmem_inst/N23 ) );
  AOI22_X1 U1122 ( .A1(n1098), .A2(\xmem_inst/mem[12][7] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][7] ), .ZN(n981) );
  AOI22_X1 U1123 ( .A1(n1099), .A2(\xmem_inst/mem[14][7] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][7] ), .ZN(n980) );
  AOI22_X1 U1124 ( .A1(n1100), .A2(\xmem_inst/mem[0][7] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][7] ), .ZN(n979) );
  AOI22_X1 U1125 ( .A1(n1101), .A2(\xmem_inst/mem[2][7] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][7] ), .ZN(n978) );
  NAND4_X1 U1126 ( .A1(n981), .A2(n980), .A3(n979), .A4(n978), .ZN(n989) );
  AOI22_X1 U1127 ( .A1(n1106), .A2(\xmem_inst/mem[4][7] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][7] ), .ZN(n982) );
  OAI21_X1 U1128 ( .B1(n1767), .B2(n1855), .A(n982), .ZN(n988) );
  NAND2_X1 U1129 ( .A1(n1779), .A2(\xmem_inst/mem[11][7] ), .ZN(n986) );
  AOI22_X1 U1130 ( .A1(n1109), .A2(\xmem_inst/mem[6][7] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][7] ), .ZN(n985) );
  NAND2_X1 U1131 ( .A1(n1773), .A2(\xmem_inst/mem[9][7] ), .ZN(n984) );
  NAND2_X1 U1132 ( .A1(n1110), .A2(\xmem_inst/mem[10][7] ), .ZN(n983) );
  NAND4_X1 U1133 ( .A1(n986), .A2(n985), .A3(n984), .A4(n983), .ZN(n987) );
  OR3_X1 U1134 ( .A1(n989), .A2(n988), .A3(n987), .ZN(\xmem_inst/N22 ) );
  AOI22_X1 U1135 ( .A1(n1098), .A2(\xmem_inst/mem[12][8] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][8] ), .ZN(n993) );
  AOI22_X1 U1136 ( .A1(n1099), .A2(\xmem_inst/mem[14][8] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][8] ), .ZN(n992) );
  AOI22_X1 U1137 ( .A1(n1100), .A2(\xmem_inst/mem[0][8] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][8] ), .ZN(n991) );
  AOI22_X1 U1138 ( .A1(n1101), .A2(\xmem_inst/mem[2][8] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][8] ), .ZN(n990) );
  NAND4_X1 U1139 ( .A1(n993), .A2(n992), .A3(n991), .A4(n990), .ZN(n1001) );
  AOI22_X1 U1140 ( .A1(n1106), .A2(\xmem_inst/mem[4][8] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][8] ), .ZN(n994) );
  OAI21_X1 U1141 ( .B1(n1767), .B2(n1856), .A(n994), .ZN(n1000) );
  NAND2_X1 U1142 ( .A1(n1779), .A2(\xmem_inst/mem[11][8] ), .ZN(n998) );
  AOI22_X1 U1143 ( .A1(n1109), .A2(\xmem_inst/mem[6][8] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][8] ), .ZN(n997) );
  NAND2_X1 U1144 ( .A1(n1773), .A2(\xmem_inst/mem[9][8] ), .ZN(n996) );
  NAND2_X1 U1145 ( .A1(n1110), .A2(\xmem_inst/mem[10][8] ), .ZN(n995) );
  NAND4_X1 U1146 ( .A1(n998), .A2(n997), .A3(n996), .A4(n995), .ZN(n999) );
  OR3_X1 U1147 ( .A1(n1001), .A2(n1000), .A3(n999), .ZN(\xmem_inst/N21 ) );
  AOI22_X1 U1148 ( .A1(n1098), .A2(\xmem_inst/mem[12][9] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][9] ), .ZN(n1005) );
  AOI22_X1 U1149 ( .A1(n1099), .A2(\xmem_inst/mem[14][9] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][9] ), .ZN(n1004) );
  AOI22_X1 U1150 ( .A1(n1100), .A2(\xmem_inst/mem[0][9] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][9] ), .ZN(n1003) );
  AOI22_X1 U1151 ( .A1(n1101), .A2(\xmem_inst/mem[2][9] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][9] ), .ZN(n1002) );
  NAND4_X1 U1152 ( .A1(n1005), .A2(n1004), .A3(n1003), .A4(n1002), .ZN(n1013)
         );
  AOI22_X1 U1153 ( .A1(n1106), .A2(\xmem_inst/mem[4][9] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][9] ), .ZN(n1006) );
  OAI21_X1 U1154 ( .B1(n1767), .B2(n1857), .A(n1006), .ZN(n1012) );
  NAND2_X1 U1155 ( .A1(n1779), .A2(\xmem_inst/mem[11][9] ), .ZN(n1010) );
  AOI22_X1 U1156 ( .A1(n1109), .A2(\xmem_inst/mem[6][9] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][9] ), .ZN(n1009) );
  NAND2_X1 U1157 ( .A1(n1773), .A2(\xmem_inst/mem[9][9] ), .ZN(n1008) );
  NAND2_X1 U1158 ( .A1(n1110), .A2(\xmem_inst/mem[10][9] ), .ZN(n1007) );
  NAND4_X1 U1159 ( .A1(n1010), .A2(n1009), .A3(n1008), .A4(n1007), .ZN(n1011)
         );
  OR3_X1 U1160 ( .A1(n1013), .A2(n1012), .A3(n1011), .ZN(\xmem_inst/N20 ) );
  AOI22_X1 U1161 ( .A1(n1098), .A2(\xmem_inst/mem[12][10] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][10] ), .ZN(n1017) );
  AOI22_X1 U1162 ( .A1(n1099), .A2(\xmem_inst/mem[14][10] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][10] ), .ZN(n1016) );
  AOI22_X1 U1163 ( .A1(n1100), .A2(\xmem_inst/mem[0][10] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][10] ), .ZN(n1015) );
  AOI22_X1 U1164 ( .A1(n1101), .A2(\xmem_inst/mem[2][10] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][10] ), .ZN(n1014) );
  NAND4_X1 U1165 ( .A1(n1017), .A2(n1016), .A3(n1015), .A4(n1014), .ZN(n1025)
         );
  AOI22_X1 U1166 ( .A1(n1106), .A2(\xmem_inst/mem[4][10] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][10] ), .ZN(n1018) );
  OAI21_X1 U1167 ( .B1(n1767), .B2(n1858), .A(n1018), .ZN(n1024) );
  NAND2_X1 U1168 ( .A1(n1779), .A2(\xmem_inst/mem[11][10] ), .ZN(n1022) );
  AOI22_X1 U1169 ( .A1(n1109), .A2(\xmem_inst/mem[6][10] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][10] ), .ZN(n1021) );
  NAND2_X1 U1170 ( .A1(n1773), .A2(\xmem_inst/mem[9][10] ), .ZN(n1020) );
  NAND2_X1 U1171 ( .A1(n1110), .A2(\xmem_inst/mem[10][10] ), .ZN(n1019) );
  NAND4_X1 U1172 ( .A1(n1022), .A2(n1021), .A3(n1020), .A4(n1019), .ZN(n1023)
         );
  OR3_X1 U1173 ( .A1(n1025), .A2(n1024), .A3(n1023), .ZN(\xmem_inst/N19 ) );
  AOI22_X1 U1174 ( .A1(n1098), .A2(\xmem_inst/mem[12][11] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][11] ), .ZN(n1029) );
  AOI22_X1 U1175 ( .A1(n1099), .A2(\xmem_inst/mem[14][11] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][11] ), .ZN(n1028) );
  AOI22_X1 U1176 ( .A1(n1100), .A2(\xmem_inst/mem[0][11] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][11] ), .ZN(n1027) );
  AOI22_X1 U1177 ( .A1(n1101), .A2(\xmem_inst/mem[2][11] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][11] ), .ZN(n1026) );
  NAND4_X1 U1178 ( .A1(n1029), .A2(n1028), .A3(n1027), .A4(n1026), .ZN(n1037)
         );
  AOI22_X1 U1179 ( .A1(n1106), .A2(\xmem_inst/mem[4][11] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][11] ), .ZN(n1030) );
  OAI21_X1 U1180 ( .B1(n1767), .B2(n1859), .A(n1030), .ZN(n1036) );
  NAND2_X1 U1181 ( .A1(n1779), .A2(\xmem_inst/mem[11][11] ), .ZN(n1034) );
  AOI22_X1 U1182 ( .A1(n1109), .A2(\xmem_inst/mem[6][11] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][11] ), .ZN(n1033) );
  NAND2_X1 U1183 ( .A1(n1773), .A2(\xmem_inst/mem[9][11] ), .ZN(n1032) );
  NAND2_X1 U1184 ( .A1(n1110), .A2(\xmem_inst/mem[10][11] ), .ZN(n1031) );
  NAND4_X1 U1185 ( .A1(n1034), .A2(n1033), .A3(n1032), .A4(n1031), .ZN(n1035)
         );
  OR3_X1 U1186 ( .A1(n1037), .A2(n1036), .A3(n1035), .ZN(\xmem_inst/N18 ) );
  AOI22_X1 U1187 ( .A1(n1098), .A2(\xmem_inst/mem[12][12] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][12] ), .ZN(n1041) );
  AOI22_X1 U1188 ( .A1(n1099), .A2(\xmem_inst/mem[14][12] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][12] ), .ZN(n1040) );
  AOI22_X1 U1189 ( .A1(n1100), .A2(\xmem_inst/mem[0][12] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][12] ), .ZN(n1039) );
  AOI22_X1 U1190 ( .A1(n1101), .A2(\xmem_inst/mem[2][12] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][12] ), .ZN(n1038) );
  NAND4_X1 U1191 ( .A1(n1041), .A2(n1040), .A3(n1039), .A4(n1038), .ZN(n1049)
         );
  AOI22_X1 U1192 ( .A1(n1106), .A2(\xmem_inst/mem[4][12] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][12] ), .ZN(n1042) );
  OAI21_X1 U1193 ( .B1(n1767), .B2(n1860), .A(n1042), .ZN(n1048) );
  NAND2_X1 U1194 ( .A1(n1779), .A2(\xmem_inst/mem[11][12] ), .ZN(n1046) );
  AOI22_X1 U1195 ( .A1(n1109), .A2(\xmem_inst/mem[6][12] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][12] ), .ZN(n1045) );
  NAND2_X1 U1196 ( .A1(n1773), .A2(\xmem_inst/mem[9][12] ), .ZN(n1044) );
  NAND2_X1 U1197 ( .A1(n1110), .A2(\xmem_inst/mem[10][12] ), .ZN(n1043) );
  NAND4_X1 U1198 ( .A1(n1046), .A2(n1045), .A3(n1044), .A4(n1043), .ZN(n1047)
         );
  OR3_X1 U1199 ( .A1(n1049), .A2(n1048), .A3(n1047), .ZN(\xmem_inst/N17 ) );
  AOI22_X1 U1200 ( .A1(n1098), .A2(\xmem_inst/mem[12][13] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][13] ), .ZN(n1053) );
  AOI22_X1 U1201 ( .A1(n1099), .A2(\xmem_inst/mem[14][13] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][13] ), .ZN(n1052) );
  AOI22_X1 U1202 ( .A1(n1100), .A2(\xmem_inst/mem[0][13] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][13] ), .ZN(n1051) );
  AOI22_X1 U1203 ( .A1(n1101), .A2(\xmem_inst/mem[2][13] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][13] ), .ZN(n1050) );
  NAND4_X1 U1204 ( .A1(n1053), .A2(n1052), .A3(n1051), .A4(n1050), .ZN(n1061)
         );
  AOI22_X1 U1205 ( .A1(n1106), .A2(\xmem_inst/mem[4][13] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][13] ), .ZN(n1054) );
  OAI21_X1 U1206 ( .B1(n1767), .B2(n1861), .A(n1054), .ZN(n1060) );
  NAND2_X1 U1207 ( .A1(n1779), .A2(\xmem_inst/mem[11][13] ), .ZN(n1058) );
  AOI22_X1 U1208 ( .A1(n1109), .A2(\xmem_inst/mem[6][13] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][13] ), .ZN(n1057) );
  NAND2_X1 U1209 ( .A1(n1773), .A2(\xmem_inst/mem[9][13] ), .ZN(n1056) );
  NAND2_X1 U1210 ( .A1(n1110), .A2(\xmem_inst/mem[10][13] ), .ZN(n1055) );
  NAND4_X1 U1211 ( .A1(n1058), .A2(n1057), .A3(n1056), .A4(n1055), .ZN(n1059)
         );
  OR3_X1 U1212 ( .A1(n1061), .A2(n1060), .A3(n1059), .ZN(\xmem_inst/N16 ) );
  AOI22_X1 U1213 ( .A1(n1098), .A2(\xmem_inst/mem[12][14] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][14] ), .ZN(n1065) );
  AOI22_X1 U1214 ( .A1(n1099), .A2(\xmem_inst/mem[14][14] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][14] ), .ZN(n1064) );
  AOI22_X1 U1215 ( .A1(n1100), .A2(\xmem_inst/mem[0][14] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][14] ), .ZN(n1063) );
  AOI22_X1 U1216 ( .A1(n1101), .A2(\xmem_inst/mem[2][14] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][14] ), .ZN(n1062) );
  NAND4_X1 U1217 ( .A1(n1065), .A2(n1064), .A3(n1063), .A4(n1062), .ZN(n1073)
         );
  AOI22_X1 U1218 ( .A1(n1106), .A2(\xmem_inst/mem[4][14] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][14] ), .ZN(n1066) );
  OAI21_X1 U1219 ( .B1(n1767), .B2(n1862), .A(n1066), .ZN(n1072) );
  NAND2_X1 U1220 ( .A1(n1779), .A2(\xmem_inst/mem[11][14] ), .ZN(n1070) );
  AOI22_X1 U1221 ( .A1(n1109), .A2(\xmem_inst/mem[6][14] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][14] ), .ZN(n1069) );
  NAND2_X1 U1222 ( .A1(n1773), .A2(\xmem_inst/mem[9][14] ), .ZN(n1068) );
  NAND2_X1 U1223 ( .A1(n1110), .A2(\xmem_inst/mem[10][14] ), .ZN(n1067) );
  NAND4_X1 U1224 ( .A1(n1070), .A2(n1069), .A3(n1068), .A4(n1067), .ZN(n1071)
         );
  OR3_X1 U1225 ( .A1(n1073), .A2(n1072), .A3(n1071), .ZN(\xmem_inst/N15 ) );
  AOI22_X1 U1226 ( .A1(n1098), .A2(\xmem_inst/mem[12][0] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][0] ), .ZN(n1077) );
  AOI22_X1 U1227 ( .A1(n1099), .A2(\xmem_inst/mem[14][0] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][0] ), .ZN(n1076) );
  AOI22_X1 U1228 ( .A1(n1100), .A2(\xmem_inst/mem[0][0] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][0] ), .ZN(n1075) );
  AOI22_X1 U1229 ( .A1(n1101), .A2(\xmem_inst/mem[2][0] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][0] ), .ZN(n1074) );
  NAND4_X1 U1230 ( .A1(n1077), .A2(n1076), .A3(n1075), .A4(n1074), .ZN(n1085)
         );
  AOI22_X1 U1231 ( .A1(n1106), .A2(\xmem_inst/mem[4][0] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][0] ), .ZN(n1078) );
  OAI21_X1 U1232 ( .B1(n1767), .B2(n1848), .A(n1078), .ZN(n1084) );
  NAND2_X1 U1233 ( .A1(n1779), .A2(\xmem_inst/mem[11][0] ), .ZN(n1082) );
  AOI22_X1 U1234 ( .A1(n1109), .A2(\xmem_inst/mem[6][0] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][0] ), .ZN(n1081) );
  NAND2_X1 U1235 ( .A1(n1773), .A2(\xmem_inst/mem[9][0] ), .ZN(n1080) );
  NAND2_X1 U1236 ( .A1(n1110), .A2(\xmem_inst/mem[10][0] ), .ZN(n1079) );
  NAND4_X1 U1237 ( .A1(n1082), .A2(n1081), .A3(n1080), .A4(n1079), .ZN(n1083)
         );
  OR3_X1 U1238 ( .A1(n1085), .A2(n1084), .A3(n1083), .ZN(\xmem_inst/N29 ) );
  AOI22_X1 U1239 ( .A1(n1098), .A2(\xmem_inst/mem[12][1] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][1] ), .ZN(n1089) );
  AOI22_X1 U1240 ( .A1(n1099), .A2(\xmem_inst/mem[14][1] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][1] ), .ZN(n1088) );
  AOI22_X1 U1241 ( .A1(n1100), .A2(\xmem_inst/mem[0][1] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][1] ), .ZN(n1087) );
  AOI22_X1 U1242 ( .A1(n1101), .A2(\xmem_inst/mem[2][1] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][1] ), .ZN(n1086) );
  NAND4_X1 U1243 ( .A1(n1089), .A2(n1088), .A3(n1087), .A4(n1086), .ZN(n1097)
         );
  AOI22_X1 U1244 ( .A1(n1106), .A2(\xmem_inst/mem[4][1] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][1] ), .ZN(n1090) );
  OAI21_X1 U1245 ( .B1(n1767), .B2(n1849), .A(n1090), .ZN(n1096) );
  NAND2_X1 U1246 ( .A1(n1779), .A2(\xmem_inst/mem[11][1] ), .ZN(n1094) );
  AOI22_X1 U1247 ( .A1(n1109), .A2(\xmem_inst/mem[6][1] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][1] ), .ZN(n1093) );
  NAND2_X1 U1248 ( .A1(n1773), .A2(\xmem_inst/mem[9][1] ), .ZN(n1092) );
  NAND2_X1 U1249 ( .A1(n1110), .A2(\xmem_inst/mem[10][1] ), .ZN(n1091) );
  NAND4_X1 U1250 ( .A1(n1094), .A2(n1093), .A3(n1092), .A4(n1091), .ZN(n1095)
         );
  OR3_X1 U1251 ( .A1(n1097), .A2(n1096), .A3(n1095), .ZN(\xmem_inst/N28 ) );
  AOI22_X1 U1252 ( .A1(n1098), .A2(\xmem_inst/mem[12][2] ), .B1(n1785), .B2(
        \xmem_inst/mem[13][2] ), .ZN(n1105) );
  AOI22_X1 U1253 ( .A1(n1099), .A2(\xmem_inst/mem[14][2] ), .B1(n1735), .B2(
        \xmem_inst/mem[15][2] ), .ZN(n1104) );
  AOI22_X1 U1254 ( .A1(n1100), .A2(\xmem_inst/mem[0][2] ), .B1(n1749), .B2(
        \xmem_inst/mem[1][2] ), .ZN(n1103) );
  AOI22_X1 U1255 ( .A1(n1101), .A2(\xmem_inst/mem[2][2] ), .B1(n1756), .B2(
        \xmem_inst/mem[3][2] ), .ZN(n1102) );
  NAND4_X1 U1256 ( .A1(n1105), .A2(n1104), .A3(n1103), .A4(n1102), .ZN(n1117)
         );
  AOI22_X1 U1257 ( .A1(n1106), .A2(\xmem_inst/mem[4][2] ), .B1(n1761), .B2(
        \xmem_inst/mem[5][2] ), .ZN(n1107) );
  OAI21_X1 U1258 ( .B1(n1767), .B2(n1850), .A(n1107), .ZN(n1116) );
  NAND2_X1 U1259 ( .A1(n1779), .A2(\xmem_inst/mem[11][2] ), .ZN(n1114) );
  AOI22_X1 U1260 ( .A1(n1109), .A2(\xmem_inst/mem[6][2] ), .B1(n1108), .B2(
        \xmem_inst/mem[8][2] ), .ZN(n1113) );
  NAND2_X1 U1261 ( .A1(n1773), .A2(\xmem_inst/mem[9][2] ), .ZN(n1112) );
  NAND2_X1 U1262 ( .A1(n1110), .A2(\xmem_inst/mem[10][2] ), .ZN(n1111) );
  NAND4_X1 U1263 ( .A1(n1114), .A2(n1113), .A3(n1112), .A4(n1111), .ZN(n1115)
         );
  OR3_X1 U1264 ( .A1(n1117), .A2(n1116), .A3(n1115), .ZN(\xmem_inst/N27 ) );
  NOR2_X1 U1265 ( .A1(n1865), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[1]) );
  NOR2_X1 U1266 ( .A1(n1843), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[8]) );
  NOR2_X1 U1267 ( .A1(n1873), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[11]) );
  NOR2_X1 U1268 ( .A1(n1867), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[6]) );
  NOR2_X1 U1269 ( .A1(n1874), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[13]) );
  NOR2_X1 U1270 ( .A1(n1866), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[2]) );
  NOR2_X1 U1271 ( .A1(n1864), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[3]) );
  NOR2_X1 U1272 ( .A1(n1871), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[5]) );
  NOR2_X1 U1273 ( .A1(n1869), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[4]) );
  NOR2_X1 U1274 ( .A1(n1846), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[12]) );
  NOR2_X1 U1275 ( .A1(n1844), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[9]) );
  NOR2_X1 U1276 ( .A1(n1872), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[7]) );
  NOR2_X1 U1277 ( .A1(n1847), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[14]) );
  NOR2_X1 U1278 ( .A1(n1868), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[0]) );
  NOR2_X1 U1279 ( .A1(n1845), .A2(\mac_unit_inst/adder_reg [15]), .ZN(
        m_data_out_y[10]) );
  NAND2_X1 U1280 ( .A1(m_ready_y), .A2(m_valid_y), .ZN(n1811) );
  INV_X1 U1281 ( .A(n1811), .ZN(n1727) );
  NOR2_X1 U1282 ( .A1(n2117), .A2(s_ready_x), .ZN(n1725) );
  INV_X1 U1283 ( .A(n1725), .ZN(n1169) );
  NOR2_X1 U1284 ( .A1(n1727), .A2(n1169), .ZN(n1119) );
  INV_X1 U1285 ( .A(reset), .ZN(n1812) );
  NAND2_X1 U1286 ( .A1(n1119), .A2(n1812), .ZN(n1814) );
  INV_X1 U1287 ( .A(n1814), .ZN(n2133) );
  INV_X1 U1288 ( .A(m_ready_y), .ZN(n1134) );
  NAND3_X1 U1289 ( .A1(n1134), .A2(m_valid_y), .A3(n1812), .ZN(n1118) );
  OAI21_X1 U1290 ( .B1(n1814), .B2(n1870), .A(n1118), .ZN(n874) );
  NAND2_X1 U1291 ( .A1(n1119), .A2(n1836), .ZN(n1124) );
  NOR2_X1 U1292 ( .A1(n1811), .A2(n1169), .ZN(n1120) );
  NOR2_X1 U1293 ( .A1(conv_done), .A2(reset), .ZN(n1736) );
  INV_X1 U1294 ( .A(n1736), .ZN(n1467) );
  OR2_X1 U1295 ( .A1(n1120), .A2(n1467), .ZN(n1125) );
  NOR2_X1 U1296 ( .A1(n1124), .A2(n1834), .ZN(n1121) );
  AOI211_X1 U1297 ( .C1(n1124), .C2(n1834), .A(n1125), .B(n1121), .ZN(n578) );
  XNOR2_X1 U1298 ( .A(n1121), .B(\fmem_inst/N12 ), .ZN(n1122) );
  NOR2_X1 U1299 ( .A1(n1122), .A2(n1125), .ZN(n579) );
  NOR2_X1 U1300 ( .A1(xmem_addr[2]), .A2(n1123), .ZN(n1131) );
  NAND2_X1 U1301 ( .A1(n1124), .A2(n1768), .ZN(n1126) );
  NAND2_X1 U1302 ( .A1(n1736), .A2(n1126), .ZN(n1745) );
  INV_X1 U1303 ( .A(n1745), .ZN(n1130) );
  NOR2_X1 U1304 ( .A1(n1126), .A2(n1125), .ZN(n1739) );
  INV_X1 U1305 ( .A(n1739), .ZN(n1738) );
  OAI21_X1 U1306 ( .B1(n1127), .B2(n1745), .A(n1738), .ZN(n1742) );
  NOR3_X1 U1307 ( .A1(n1467), .A2(n1811), .A3(n1169), .ZN(n1743) );
  AOI22_X1 U1308 ( .A1(xmem_addr[2]), .A2(n1742), .B1(n1743), .B2(
        \ctrl_conv_output_inst/cnt_conv [2]), .ZN(n1128) );
  INV_X1 U1309 ( .A(n1128), .ZN(n1129) );
  AOI21_X1 U1310 ( .B1(n1131), .B2(n1130), .A(n1129), .ZN(n1132) );
  INV_X1 U1311 ( .A(n1132), .ZN(n870) );
  AND2_X1 U1312 ( .A1(\ctrl_conv_output_inst/conv_start_accum ), .A2(n1812), 
        .ZN(n1462) );
  AND2_X1 U1313 ( .A1(n1462), .A2(m_valid_y), .ZN(n1133) );
  NAND2_X1 U1314 ( .A1(n1134), .A2(n1133), .ZN(n1591) );
  NOR2_X1 U1315 ( .A1(\mac_unit_inst/adder_reg [2]), .A2(
        \mac_unit_inst/x_mult_f_reg [2]), .ZN(n1492) );
  NOR2_X1 U1316 ( .A1(\mac_unit_inst/adder_reg [3]), .A2(
        \mac_unit_inst/x_mult_f_reg [3]), .ZN(n1494) );
  NOR2_X1 U1317 ( .A1(n1492), .A2(n1494), .ZN(n1136) );
  NOR2_X1 U1318 ( .A1(\mac_unit_inst/adder_reg [1]), .A2(
        \mac_unit_inst/x_mult_f_reg [1]), .ZN(n1479) );
  NAND2_X1 U1319 ( .A1(\mac_unit_inst/adder_reg [0]), .A2(
        \mac_unit_inst/x_mult_f_reg [0]), .ZN(n1482) );
  NAND2_X1 U1320 ( .A1(\mac_unit_inst/adder_reg [1]), .A2(
        \mac_unit_inst/x_mult_f_reg [1]), .ZN(n1480) );
  OAI21_X1 U1321 ( .B1(n1479), .B2(n1482), .A(n1480), .ZN(n1486) );
  NAND2_X1 U1322 ( .A1(\mac_unit_inst/adder_reg [2]), .A2(
        \mac_unit_inst/x_mult_f_reg [2]), .ZN(n1491) );
  NAND2_X1 U1323 ( .A1(\mac_unit_inst/adder_reg [3]), .A2(
        \mac_unit_inst/x_mult_f_reg [3]), .ZN(n1495) );
  OAI21_X1 U1324 ( .B1(n1494), .B2(n1491), .A(n1495), .ZN(n1135) );
  AOI21_X1 U1325 ( .B1(n1136), .B2(n1486), .A(n1135), .ZN(n1501) );
  NOR2_X1 U1326 ( .A1(\mac_unit_inst/adder_reg [4]), .A2(
        \mac_unit_inst/x_mult_f_reg [4]), .ZN(n1502) );
  NOR2_X1 U1327 ( .A1(\mac_unit_inst/adder_reg [5]), .A2(
        \mac_unit_inst/x_mult_f_reg [5]), .ZN(n1509) );
  NOR2_X1 U1328 ( .A1(n1502), .A2(n1509), .ZN(n1517) );
  NOR2_X1 U1329 ( .A1(\mac_unit_inst/adder_reg [6]), .A2(
        \mac_unit_inst/x_mult_f_reg [6]), .ZN(n1524) );
  NOR2_X1 U1330 ( .A1(\mac_unit_inst/adder_reg [7]), .A2(
        \mac_unit_inst/x_mult_f_reg [7]), .ZN(n1526) );
  NOR2_X1 U1331 ( .A1(n1524), .A2(n1526), .ZN(n1138) );
  NAND2_X1 U1332 ( .A1(n1517), .A2(n1138), .ZN(n1140) );
  NAND2_X1 U1333 ( .A1(\mac_unit_inst/adder_reg [4]), .A2(
        \mac_unit_inst/x_mult_f_reg [4]), .ZN(n1506) );
  NAND2_X1 U1334 ( .A1(\mac_unit_inst/adder_reg [5]), .A2(
        \mac_unit_inst/x_mult_f_reg [5]), .ZN(n1510) );
  OAI21_X1 U1335 ( .B1(n1509), .B2(n1506), .A(n1510), .ZN(n1516) );
  NAND2_X1 U1336 ( .A1(\mac_unit_inst/adder_reg [6]), .A2(
        \mac_unit_inst/x_mult_f_reg [6]), .ZN(n1523) );
  NAND2_X1 U1337 ( .A1(\mac_unit_inst/adder_reg [7]), .A2(
        \mac_unit_inst/x_mult_f_reg [7]), .ZN(n1527) );
  OAI21_X1 U1338 ( .B1(n1526), .B2(n1523), .A(n1527), .ZN(n1137) );
  AOI21_X1 U1339 ( .B1(n1138), .B2(n1516), .A(n1137), .ZN(n1139) );
  OAI21_X1 U1340 ( .B1(n1501), .B2(n1140), .A(n1139), .ZN(n1533) );
  NOR2_X1 U1341 ( .A1(\mac_unit_inst/adder_reg [8]), .A2(
        \mac_unit_inst/x_mult_f_reg [8]), .ZN(n1582) );
  NOR2_X1 U1342 ( .A1(\mac_unit_inst/adder_reg [9]), .A2(
        \mac_unit_inst/x_mult_f_reg [9]), .ZN(n1534) );
  NOR2_X1 U1343 ( .A1(n1582), .A2(n1534), .ZN(n1541) );
  NOR2_X1 U1344 ( .A1(\mac_unit_inst/adder_reg [10]), .A2(
        \mac_unit_inst/x_mult_f_reg [10]), .ZN(n1545) );
  NOR2_X1 U1345 ( .A1(\mac_unit_inst/adder_reg [11]), .A2(
        \mac_unit_inst/x_mult_f_reg [11]), .ZN(n1553) );
  NOR2_X1 U1346 ( .A1(n1545), .A2(n1553), .ZN(n1143) );
  NAND2_X1 U1347 ( .A1(n1541), .A2(n1143), .ZN(n1153) );
  INV_X1 U1348 ( .A(n1153), .ZN(n1141) );
  NAND2_X1 U1349 ( .A1(n1533), .A2(n1141), .ZN(n1144) );
  NAND2_X1 U1350 ( .A1(\mac_unit_inst/adder_reg [8]), .A2(
        \mac_unit_inst/x_mult_f_reg [8]), .ZN(n1583) );
  NAND2_X1 U1351 ( .A1(\mac_unit_inst/adder_reg [9]), .A2(
        \mac_unit_inst/x_mult_f_reg [9]), .ZN(n1535) );
  OAI21_X1 U1352 ( .B1(n1534), .B2(n1583), .A(n1535), .ZN(n1542) );
  NAND2_X1 U1353 ( .A1(\mac_unit_inst/adder_reg [10]), .A2(
        \mac_unit_inst/x_mult_f_reg [10]), .ZN(n1549) );
  NAND2_X1 U1354 ( .A1(\mac_unit_inst/adder_reg [11]), .A2(
        \mac_unit_inst/x_mult_f_reg [11]), .ZN(n1554) );
  OAI21_X1 U1355 ( .B1(n1553), .B2(n1549), .A(n1554), .ZN(n1142) );
  AOI21_X1 U1356 ( .B1(n1143), .B2(n1542), .A(n1142), .ZN(n1160) );
  NAND2_X1 U1357 ( .A1(n1144), .A2(n1160), .ZN(n1568) );
  NOR2_X1 U1358 ( .A1(\mac_unit_inst/adder_reg [12]), .A2(
        \mac_unit_inst/x_mult_f_reg [12]), .ZN(n1560) );
  NOR2_X1 U1359 ( .A1(\mac_unit_inst/adder_reg [13]), .A2(
        \mac_unit_inst/x_mult_f_reg [13]), .ZN(n1569) );
  NOR2_X1 U1360 ( .A1(n1560), .A2(n1569), .ZN(n1152) );
  NAND2_X1 U1361 ( .A1(n1568), .A2(n1152), .ZN(n1146) );
  NAND2_X1 U1362 ( .A1(\mac_unit_inst/adder_reg [12]), .A2(
        \mac_unit_inst/x_mult_f_reg [12]), .ZN(n1565) );
  NAND2_X1 U1363 ( .A1(\mac_unit_inst/adder_reg [13]), .A2(
        \mac_unit_inst/x_mult_f_reg [13]), .ZN(n1570) );
  OAI21_X1 U1364 ( .B1(n1569), .B2(n1565), .A(n1570), .ZN(n1157) );
  INV_X1 U1365 ( .A(n1157), .ZN(n1145) );
  NAND2_X1 U1366 ( .A1(n1146), .A2(n1145), .ZN(n1579) );
  NOR2_X1 U1367 ( .A1(\mac_unit_inst/adder_reg [14]), .A2(
        \mac_unit_inst/x_mult_f_reg [14]), .ZN(n1151) );
  INV_X1 U1368 ( .A(n1151), .ZN(n1577) );
  NAND2_X1 U1369 ( .A1(\mac_unit_inst/adder_reg [14]), .A2(
        \mac_unit_inst/x_mult_f_reg [14]), .ZN(n1576) );
  INV_X1 U1370 ( .A(n1576), .ZN(n1147) );
  AOI21_X1 U1371 ( .B1(n1579), .B2(n1577), .A(n1147), .ZN(n1150) );
  NOR2_X1 U1372 ( .A1(n1839), .A2(n1822), .ZN(n1155) );
  INV_X1 U1373 ( .A(n1155), .ZN(n1148) );
  NAND2_X1 U1374 ( .A1(n1839), .A2(n1822), .ZN(n1154) );
  NAND2_X1 U1375 ( .A1(n1148), .A2(n1154), .ZN(n1149) );
  XOR2_X1 U1376 ( .A(n1150), .B(n1149), .Z(n1167) );
  NOR2_X1 U1377 ( .A1(n1155), .A2(n1151), .ZN(n1158) );
  NAND2_X1 U1378 ( .A1(n1158), .A2(n1152), .ZN(n1161) );
  NOR2_X1 U1379 ( .A1(n1161), .A2(n1153), .ZN(n1163) );
  OAI21_X1 U1380 ( .B1(n1155), .B2(n1576), .A(n1154), .ZN(n1156) );
  AOI21_X1 U1381 ( .B1(n1158), .B2(n1157), .A(n1156), .ZN(n1159) );
  OAI21_X1 U1382 ( .B1(n1161), .B2(n1160), .A(n1159), .ZN(n1162) );
  AOI21_X1 U1383 ( .B1(n1163), .B2(n1533), .A(n1162), .ZN(n1164) );
  INV_X1 U1384 ( .A(n1164), .ZN(n1165) );
  NOR2_X1 U1385 ( .A1(n1167), .A2(n1165), .ZN(n1473) );
  INV_X1 U1386 ( .A(n1477), .ZN(n1166) );
  AND2_X1 U1387 ( .A1(n1462), .A2(n2035), .ZN(n1476) );
  OAI211_X1 U1388 ( .C1(n1473), .C2(n1167), .A(n1166), .B(n1476), .ZN(n1168)
         );
  OAI21_X1 U1389 ( .B1(n1839), .B2(n1591), .A(n1168), .ZN(n580) );
  NAND3_X1 U1390 ( .A1(n1811), .A2(n1462), .A3(n1169), .ZN(n1723) );
  OR2_X1 U1391 ( .A1(n1819), .A2(n1818), .ZN(n1213) );
  NAND2_X1 U1392 ( .A1(fmem_data[4]), .A2(xmem_data[13]), .ZN(n1231) );
  INV_X1 U1393 ( .A(fmem_data[4]), .ZN(n1326) );
  NOR2_X1 U1394 ( .A1(n1326), .A2(n906), .ZN(n1182) );
  AND2_X1 U1395 ( .A1(fmem_data[4]), .A2(xmem_data[11]), .ZN(n1181) );
  XNOR2_X1 U1396 ( .A(n1208), .B(n1209), .ZN(n1175) );
  AND2_X1 U1397 ( .A1(n1821), .A2(xmem_data[9]), .ZN(n1307) );
  OR2_X1 U1398 ( .A1(n1820), .A2(n1827), .ZN(n1200) );
  OR2_X1 U1399 ( .A1(n881), .A2(n1826), .ZN(n1251) );
  INV_X1 U1400 ( .A(n1251), .ZN(n1171) );
  OR2_X1 U1401 ( .A1(n1819), .A2(n909), .ZN(n1183) );
  INV_X1 U1402 ( .A(n1183), .ZN(n1170) );
  NAND2_X1 U1403 ( .A1(n1171), .A2(n1170), .ZN(n1172) );
  NAND2_X1 U1404 ( .A1(n1185), .A2(n1172), .ZN(n1174) );
  NAND2_X1 U1405 ( .A1(n1183), .A2(n1251), .ZN(n1173) );
  NAND2_X1 U1406 ( .A1(n1174), .A2(n1173), .ZN(n1207) );
  XNOR2_X1 U1407 ( .A(n1175), .B(n1207), .ZN(n1411) );
  NOR2_X1 U1408 ( .A1(n1820), .A2(n1818), .ZN(n1191) );
  NOR2_X1 U1409 ( .A1(n1283), .A2(n907), .ZN(n1190) );
  NOR2_X1 U1410 ( .A1(n881), .A2(n1817), .ZN(n1228) );
  OR2_X1 U1411 ( .A1(n1819), .A2(n1815), .ZN(n1202) );
  INV_X1 U1412 ( .A(n1202), .ZN(n1177) );
  INV_X1 U1413 ( .A(n1201), .ZN(n1176) );
  NAND2_X1 U1414 ( .A1(n1204), .A2(n1178), .ZN(n1180) );
  NAND2_X1 U1415 ( .A1(n1202), .A2(n1201), .ZN(n1179) );
  NAND2_X1 U1416 ( .A1(n1180), .A2(n1179), .ZN(n1220) );
  FA_X1 U1417 ( .A(n1182), .B(n1181), .CI(n1298), .CO(n1209), .S(n1219) );
  XNOR2_X1 U1418 ( .A(n1251), .B(n1183), .ZN(n1184) );
  XNOR2_X1 U1419 ( .A(n1185), .B(n1184), .ZN(n1218) );
  INV_X1 U1420 ( .A(n1412), .ZN(n1186) );
  XNOR2_X1 U1421 ( .A(n1411), .B(n1186), .ZN(n1256) );
  NOR2_X1 U1422 ( .A1(n1820), .A2(n1815), .ZN(n1281) );
  OR2_X1 U1423 ( .A1(n1819), .A2(n911), .ZN(n1274) );
  NOR2_X2 U1424 ( .A1(n882), .A2(n908), .ZN(n1355) );
  NAND2_X1 U1425 ( .A1(n1276), .A2(n1187), .ZN(n1189) );
  NAND2_X1 U1426 ( .A1(n1189), .A2(n1188), .ZN(n1289) );
  FA_X1 U1427 ( .A(n1191), .B(n1190), .CI(n1228), .CO(n1204), .S(n1288) );
  NOR2_X1 U1428 ( .A1(n1820), .A2(n909), .ZN(n1273) );
  NOR2_X1 U1429 ( .A1(n1817), .A2(n1283), .ZN(n1272) );
  NOR2_X2 U1430 ( .A1(n881), .A2(n1815), .ZN(n1367) );
  OR2_X1 U1431 ( .A1(n1819), .A2(n908), .ZN(n1197) );
  XNOR2_X1 U1432 ( .A(n1367), .B(n1197), .ZN(n1192) );
  XNOR2_X1 U1433 ( .A(n1196), .B(n1192), .ZN(n1287) );
  INV_X1 U1434 ( .A(n1367), .ZN(n1194) );
  INV_X1 U1435 ( .A(n1197), .ZN(n1193) );
  NAND2_X1 U1436 ( .A1(n1194), .A2(n1193), .ZN(n1195) );
  NAND2_X1 U1437 ( .A1(n1196), .A2(n1195), .ZN(n1199) );
  NAND2_X1 U1438 ( .A1(n1367), .A2(n1197), .ZN(n1198) );
  NAND2_X1 U1439 ( .A1(n1199), .A2(n1198), .ZN(n1221) );
  FA_X1 U1440 ( .A(n1307), .B(n1250), .CI(n1200), .CO(n1185), .S(n1223) );
  XNOR2_X1 U1441 ( .A(n1202), .B(n1201), .ZN(n1203) );
  XNOR2_X1 U1442 ( .A(n1204), .B(n1203), .ZN(n1222) );
  OAI21_X1 U1443 ( .B1(n1221), .B2(n1223), .A(n1222), .ZN(n1206) );
  NAND2_X1 U1444 ( .A1(n1223), .A2(n1221), .ZN(n1205) );
  NAND2_X1 U1445 ( .A1(n1206), .A2(n1205), .ZN(n1414) );
  OAI21_X1 U1446 ( .B1(n1209), .B2(n1208), .A(n1207), .ZN(n1212) );
  BUF_X1 U1447 ( .A(n1208), .Z(n1210) );
  NAND2_X1 U1448 ( .A1(n1210), .A2(n1209), .ZN(n1211) );
  NAND2_X1 U1449 ( .A1(n1212), .A2(n1211), .ZN(n1433) );
  INV_X1 U1450 ( .A(n1433), .ZN(n1215) );
  FA_X1 U1451 ( .A(n1213), .B(n1231), .CI(n886), .CO(n1422), .S(n1208) );
  INV_X1 U1452 ( .A(fmem_data[15]), .ZN(n1350) );
  OR2_X1 U1453 ( .A1(n1350), .A2(n1827), .ZN(n1421) );
  NOR2_X1 U1454 ( .A1(n1820), .A2(n907), .ZN(n1232) );
  XNOR2_X1 U1455 ( .A(n1214), .B(n1215), .ZN(n1257) );
  OAI21_X1 U1456 ( .B1(n1256), .B2(n910), .A(n1257), .ZN(n1216) );
  INV_X1 U1457 ( .A(n1216), .ZN(n1597) );
  INV_X1 U1458 ( .A(n1414), .ZN(n1217) );
  XNOR2_X1 U1459 ( .A(n1217), .B(n1415), .ZN(n1225) );
  FA_X1 U1460 ( .A(n1220), .B(n1219), .CI(n1218), .CO(n1412), .S(n1426) );
  NOR2_X1 U1461 ( .A1(n1225), .A2(n1426), .ZN(n1595) );
  INV_X1 U1462 ( .A(n1415), .ZN(n1416) );
  NAND2_X1 U1463 ( .A1(n1417), .A2(n1416), .ZN(n1429) );
  NAND2_X1 U1464 ( .A1(n1225), .A2(n1426), .ZN(n1226) );
  OAI21_X1 U1465 ( .B1(n1595), .B2(n1429), .A(n1226), .ZN(n1227) );
  NAND2_X1 U1466 ( .A1(n1597), .A2(n1227), .ZN(n1265) );
  OR2_X1 U1467 ( .A1(n1350), .A2(n1817), .ZN(n1241) );
  INV_X1 U1468 ( .A(n1250), .ZN(n1240) );
  INV_X1 U1469 ( .A(n1231), .ZN(n1233) );
  OAI21_X1 U1470 ( .B1(n1228), .B2(n1233), .A(n1234), .ZN(n1230) );
  NOR2_X1 U1471 ( .A1(n882), .A2(n1817), .ZN(n1235) );
  NAND2_X1 U1472 ( .A1(n1235), .A2(n1233), .ZN(n1229) );
  NAND2_X1 U1473 ( .A1(n1230), .A2(n1229), .ZN(n1239) );
  FA_X1 U1474 ( .A(n1271), .B(n1232), .CI(n895), .CO(n1246), .S(n1420) );
  OR2_X1 U1475 ( .A1(n1350), .A2(n906), .ZN(n1244) );
  XNOR2_X1 U1476 ( .A(n1234), .B(n1233), .ZN(n1236) );
  XNOR2_X1 U1477 ( .A(n1236), .B(n1235), .ZN(n1247) );
  OAI21_X1 U1478 ( .B1(n1246), .B2(n1244), .A(n1247), .ZN(n1238) );
  XOR2_X1 U1479 ( .A(n1442), .B(n1441), .Z(n1243) );
  FA_X1 U1480 ( .A(n1241), .B(n1240), .CI(n1239), .CO(n1444), .S(n1442) );
  OR2_X1 U1481 ( .A1(n1350), .A2(n907), .ZN(n1249) );
  NAND2_X1 U1482 ( .A1(n1243), .A2(n1242), .ZN(n1255) );
  FA_X1 U1483 ( .A(n1422), .B(n1421), .CI(n1420), .CO(n1440), .S(n1214) );
  INV_X1 U1484 ( .A(n1244), .ZN(n1245) );
  XNOR2_X1 U1485 ( .A(n1246), .B(n1245), .ZN(n1248) );
  XNOR2_X1 U1486 ( .A(n1248), .B(n1247), .ZN(n1419) );
  XNOR2_X1 U1487 ( .A(n1440), .B(n1419), .ZN(n1253) );
  FA_X1 U1488 ( .A(n1251), .B(n1250), .CI(n1249), .CO(n1451), .S(n1443) );
  NOR2_X1 U1489 ( .A1(n1350), .A2(n1826), .ZN(n1450) );
  HA_X1 U1490 ( .A(n1451), .B(n1450), .S(n1252) );
  NAND2_X1 U1491 ( .A1(n1253), .A2(n1252), .ZN(n1254) );
  INV_X1 U1492 ( .A(n1598), .ZN(n1263) );
  NAND2_X1 U1493 ( .A1(n1256), .A2(n910), .ZN(n1261) );
  INV_X1 U1494 ( .A(n1257), .ZN(n1260) );
  AND2_X1 U1495 ( .A1(n1411), .A2(n903), .ZN(n1258) );
  NAND2_X1 U1496 ( .A1(n1258), .A2(n1257), .ZN(n1259) );
  OAI21_X1 U1497 ( .B1(n1261), .B2(n1260), .A(n1259), .ZN(n1262) );
  NAND2_X1 U1498 ( .A1(n1263), .A2(n1262), .ZN(n1264) );
  OAI21_X1 U1499 ( .B1(n1265), .B2(n1598), .A(n1264), .ZN(n1593) );
  INV_X1 U1500 ( .A(n892), .ZN(n1465) );
  NOR2_X1 U1501 ( .A1(n1820), .A2(n908), .ZN(n1297) );
  BUF_X2 U1502 ( .A(n1823), .Z(n1605) );
  NOR2_X1 U1503 ( .A1(n1605), .A2(n1827), .ZN(n1296) );
  OR2_X1 U1504 ( .A1(n1819), .A2(n1825), .ZN(n1277) );
  INV_X1 U1505 ( .A(n1277), .ZN(n1267) );
  INV_X1 U1506 ( .A(n1354), .ZN(n1266) );
  NAND2_X1 U1507 ( .A1(n1267), .A2(n1266), .ZN(n1268) );
  NAND2_X1 U1508 ( .A1(n1279), .A2(n1268), .ZN(n1270) );
  NAND2_X1 U1509 ( .A1(n1277), .A2(n1354), .ZN(n1269) );
  NAND2_X1 U1510 ( .A1(n1270), .A2(n1269), .ZN(n1292) );
  FA_X1 U1511 ( .A(n1273), .B(n1272), .CI(n1271), .CO(n1196), .S(n1291) );
  XNOR2_X1 U1512 ( .A(n1355), .B(n1274), .ZN(n1275) );
  XNOR2_X1 U1513 ( .A(n1276), .B(n1275), .ZN(n1290) );
  XNOR2_X1 U1514 ( .A(n1277), .B(n1354), .ZN(n1278) );
  XNOR2_X1 U1515 ( .A(n1279), .B(n1278), .ZN(n1317) );
  NOR2_X1 U1516 ( .A1(n1283), .A2(n1818), .ZN(n1309) );
  AND2_X1 U1517 ( .A1(fmem_data[4]), .A2(xmem_data[6]), .ZN(n1308) );
  OR2_X1 U1518 ( .A1(n1819), .A2(n1829), .ZN(n1299) );
  NOR2_X1 U1519 ( .A1(n882), .A2(n1825), .ZN(n1331) );
  OR2_X1 U1520 ( .A1(n1299), .A2(n1331), .ZN(n1284) );
  NAND2_X1 U1521 ( .A1(n1331), .A2(n1299), .ZN(n1285) );
  NAND2_X1 U1522 ( .A1(n1286), .A2(n1285), .ZN(n1315) );
  NOR2_X1 U1523 ( .A1(n1396), .A2(n1395), .ZN(n1700) );
  FA_X1 U1524 ( .A(n1289), .B(n1288), .CI(n1287), .CO(n1415), .S(n1398) );
  FA_X1 U1525 ( .A(n1292), .B(n1291), .CI(n1290), .CO(n1397), .S(n1396) );
  NOR2_X1 U1526 ( .A1(n1398), .A2(n1397), .ZN(n1714) );
  NOR2_X1 U1527 ( .A1(n1700), .A2(n1714), .ZN(n1400) );
  NOR2_X1 U1528 ( .A1(n1605), .A2(n909), .ZN(n1369) );
  NOR2_X1 U1529 ( .A1(n1820), .A2(n1825), .ZN(n1368) );
  OR2_X1 U1530 ( .A1(n1819), .A2(n1832), .ZN(n1310) );
  NOR2_X2 U1531 ( .A1(n882), .A2(n1829), .ZN(n1333) );
  INV_X1 U1532 ( .A(n1333), .ZN(n1293) );
  NAND2_X1 U1533 ( .A1(n1294), .A2(n1293), .ZN(n1295) );
  NAND2_X1 U1534 ( .A1(n1312), .A2(n1295), .ZN(n1319) );
  FA_X1 U1535 ( .A(n1297), .B(n1298), .CI(n1296), .CO(n1279), .S(n1323) );
  XNOR2_X1 U1536 ( .A(n1320), .B(n1323), .ZN(n1302) );
  XNOR2_X1 U1537 ( .A(n1331), .B(n1299), .ZN(n1300) );
  XNOR2_X1 U1538 ( .A(n1302), .B(n1322), .ZN(n1392) );
  INV_X1 U1539 ( .A(n1816), .ZN(n1339) );
  NOR2_X1 U1540 ( .A1(n1339), .A2(n1815), .ZN(n1357) );
  NOR2_X1 U1541 ( .A1(n1820), .A2(n1829), .ZN(n1356) );
  OR2_X1 U1542 ( .A1(n1819), .A2(n1831), .ZN(n1373) );
  FA_X1 U1543 ( .A(n1309), .B(n1308), .CI(n1307), .CO(n1301), .S(n1380) );
  XNOR2_X1 U1544 ( .A(n1333), .B(n1310), .ZN(n1311) );
  XNOR2_X1 U1545 ( .A(n1312), .B(n1311), .ZN(n1381) );
  NOR2_X1 U1546 ( .A1(n1391), .A2(n1392), .ZN(n1682) );
  FA_X1 U1547 ( .A(n1317), .B(n1316), .CI(n1315), .CO(n1395), .S(n1394) );
  NAND2_X1 U1548 ( .A1(n1319), .A2(n1318), .ZN(n1320) );
  NAND2_X1 U1549 ( .A1(n1325), .A2(n1324), .ZN(n1393) );
  NOR2_X1 U1550 ( .A1(n1682), .A2(n898), .ZN(n1697) );
  NAND2_X1 U1551 ( .A1(n1400), .A2(n1697), .ZN(n1409) );
  NOR2_X1 U1552 ( .A1(n1605), .A2(n911), .ZN(n1332) );
  INV_X1 U1553 ( .A(n881), .ZN(n1338) );
  NAND2_X1 U1554 ( .A1(n1338), .A2(xmem_data[0]), .ZN(n1327) );
  NOR2_X1 U1555 ( .A1(n1326), .A2(n1831), .ZN(n1358) );
  XNOR2_X1 U1556 ( .A(n1327), .B(n1358), .ZN(n1330) );
  AND2_X1 U1557 ( .A1(n884), .A2(n1358), .ZN(n1328) );
  AND2_X1 U1558 ( .A1(n1816), .A2(xmem_data[7]), .ZN(n1351) );
  NOR2_X1 U1559 ( .A1(n1820), .A2(n1832), .ZN(n1352) );
  XNOR2_X1 U1560 ( .A(n1351), .B(n1352), .ZN(n1361) );
  NOR2_X1 U1561 ( .A1(n882), .A2(n1830), .ZN(n1612) );
  OR2_X1 U1562 ( .A1(n1350), .A2(n1824), .ZN(n1353) );
  FA_X1 U1563 ( .A(n1332), .B(n1331), .CI(n1330), .CO(n1360), .S(n1347) );
  NOR2_X1 U1564 ( .A1(n1339), .A2(n1825), .ZN(n1335) );
  NOR2_X1 U1565 ( .A1(n1820), .A2(n1830), .ZN(n1334) );
  NOR2_X1 U1566 ( .A1(n1347), .A2(n1346), .ZN(n1642) );
  FA_X1 U1567 ( .A(n1334), .B(n1335), .CI(n1333), .CO(n1346), .S(n1345) );
  NOR2_X1 U1568 ( .A1(n1326), .A2(n1824), .ZN(n1336) );
  INV_X1 U1569 ( .A(n1374), .ZN(n1337) );
  XNOR2_X1 U1570 ( .A(n1337), .B(n1336), .ZN(n1343) );
  NOR2_X1 U1571 ( .A1(n1339), .A2(n1829), .ZN(n1342) );
  NOR2_X1 U1572 ( .A1(n1343), .A2(n1342), .ZN(n1627) );
  NOR2_X1 U1573 ( .A1(n1605), .A2(n1831), .ZN(n1613) );
  NAND2_X1 U1574 ( .A1(n1613), .A2(n1612), .ZN(n1614) );
  NOR2_X1 U1575 ( .A1(n1605), .A2(n1830), .ZN(n1608) );
  NAND3_X1 U1576 ( .A1(n1338), .A2(xmem_data[0]), .A3(n1608), .ZN(n1616) );
  NAND2_X1 U1577 ( .A1(n1614), .A2(n1616), .ZN(n1624) );
  NOR2_X1 U1578 ( .A1(n1339), .A2(n1832), .ZN(n1340) );
  NOR2_X1 U1579 ( .A1(n881), .A2(n1831), .ZN(n1371) );
  OR2_X1 U1580 ( .A1(n1340), .A2(n1371), .ZN(n1622) );
  NAND2_X1 U1581 ( .A1(n1340), .A2(n1371), .ZN(n1621) );
  INV_X1 U1582 ( .A(n1621), .ZN(n1341) );
  AOI21_X1 U1583 ( .B1(n1624), .B2(n1622), .A(n1341), .ZN(n1630) );
  NAND2_X1 U1584 ( .A1(n1343), .A2(n1342), .ZN(n1628) );
  OAI21_X1 U1585 ( .B1(n1627), .B2(n1630), .A(n1628), .ZN(n1637) );
  AOI21_X1 U1586 ( .B1(n1636), .B2(n885), .A(n1634), .ZN(n1641) );
  NAND2_X1 U1587 ( .A1(n1347), .A2(n1346), .ZN(n1643) );
  OAI21_X1 U1588 ( .B1(n1642), .B2(n894), .A(n1643), .ZN(n1651) );
  AND2_X1 U1589 ( .A1(n1349), .A2(n1348), .ZN(n1648) );
  AOI21_X1 U1590 ( .B1(n1649), .B2(n1651), .A(n1648), .ZN(n1656) );
  OR2_X1 U1591 ( .A1(n1350), .A2(n1830), .ZN(n1372) );
  OR2_X1 U1592 ( .A1(n1352), .A2(n1351), .ZN(n1370) );
  FA_X1 U1593 ( .A(n1354), .B(n1612), .CI(n1353), .CO(n1378), .S(n1348) );
  FA_X1 U1594 ( .A(n1357), .B(n1356), .CI(n1355), .CO(n1376), .S(n1377) );
  AND2_X1 U1595 ( .A1(n884), .A2(n1358), .ZN(n1362) );
  NOR2_X1 U1596 ( .A1(n1366), .A2(n1365), .ZN(n1657) );
  NAND2_X1 U1597 ( .A1(n1366), .A2(n1365), .ZN(n1658) );
  OAI21_X1 U1598 ( .B1(n1656), .B2(n1657), .A(n1658), .ZN(n1666) );
  FA_X1 U1599 ( .A(n1369), .B(n1368), .CI(n1367), .CO(n1312), .S(n1386) );
  FA_X1 U1600 ( .A(n1372), .B(n1371), .CI(n1370), .CO(n1385), .S(n1379) );
  XNOR2_X1 U1601 ( .A(n1374), .B(n1373), .ZN(n1375) );
  XNOR2_X1 U1602 ( .A(n1376), .B(n1375), .ZN(n1384) );
  FA_X1 U1603 ( .A(n1377), .B(n1378), .CI(n1379), .CO(n1387), .S(n1366) );
  NOR2_X1 U1604 ( .A1(n1388), .A2(n1387), .ZN(n1671) );
  XNOR2_X1 U1605 ( .A(n1381), .B(n1380), .ZN(n1383) );
  XNOR2_X1 U1606 ( .A(n1383), .B(n1382), .ZN(n1390) );
  FA_X1 U1607 ( .A(n1386), .B(n1385), .CI(n1384), .CO(n1389), .S(n1388) );
  NOR2_X1 U1608 ( .A1(n1390), .A2(n1389), .ZN(n1673) );
  NOR2_X1 U1609 ( .A1(n1671), .A2(n1673), .ZN(n1407) );
  NAND2_X1 U1610 ( .A1(n1388), .A2(n1387), .ZN(n1670) );
  NAND2_X1 U1611 ( .A1(n1390), .A2(n1389), .ZN(n1674) );
  OAI21_X1 U1612 ( .B1(n1673), .B2(n1670), .A(n1674), .ZN(n1406) );
  AOI21_X1 U1613 ( .B1(n1666), .B2(n1407), .A(n1406), .ZN(n1681) );
  NAND2_X1 U1614 ( .A1(n1392), .A2(n1391), .ZN(n1683) );
  NAND2_X1 U1615 ( .A1(n1394), .A2(n1393), .ZN(n1690) );
  OAI21_X1 U1616 ( .B1(n1689), .B2(n1683), .A(n1690), .ZN(n1698) );
  NAND2_X1 U1617 ( .A1(n1396), .A2(n1395), .ZN(n1709) );
  NAND2_X1 U1618 ( .A1(n1398), .A2(n1397), .ZN(n1715) );
  OAI21_X1 U1619 ( .B1(n899), .B2(n1709), .A(n1715), .ZN(n1399) );
  AOI21_X1 U1620 ( .B1(n1400), .B2(n1698), .A(n1399), .ZN(n1408) );
  OAI21_X1 U1621 ( .B1(n1409), .B2(n1681), .A(n1408), .ZN(n1405) );
  INV_X1 U1622 ( .A(n1416), .ZN(n1401) );
  OR2_X1 U1623 ( .A1(n1417), .A2(n1401), .ZN(n1403) );
  NAND2_X1 U1624 ( .A1(n1417), .A2(n1401), .ZN(n1402) );
  NAND2_X1 U1625 ( .A1(n1403), .A2(n1402), .ZN(n1404) );
  XNOR2_X1 U1626 ( .A(n1405), .B(n1404), .ZN(n1464) );
  AOI21_X1 U1627 ( .B1(n1666), .B2(n1407), .A(n1406), .ZN(n1410) );
  OAI21_X1 U1628 ( .B1(n1410), .B2(n1409), .A(n1408), .ZN(n1602) );
  XNOR2_X1 U1629 ( .A(n1411), .B(n903), .ZN(n1432) );
  OR2_X1 U1630 ( .A1(n1415), .A2(n1414), .ZN(n1431) );
  NOR2_X1 U1631 ( .A1(n1432), .A2(n1431), .ZN(n1413) );
  NOR2_X1 U1632 ( .A1(n1413), .A2(n880), .ZN(n1438) );
  XNOR2_X1 U1633 ( .A(n1415), .B(n1414), .ZN(n1427) );
  NOR2_X1 U1634 ( .A1(n1426), .A2(n1427), .ZN(n1430) );
  NOR2_X1 U1635 ( .A1(n1417), .A2(n1416), .ZN(n1594) );
  NOR2_X1 U1636 ( .A1(n1430), .A2(n1594), .ZN(n1418) );
  NAND2_X1 U1637 ( .A1(n1438), .A2(n1418), .ZN(n1424) );
  OR2_X1 U1638 ( .A1(n1442), .A2(n1441), .ZN(n1446) );
  INV_X1 U1639 ( .A(n1419), .ZN(n1439) );
  NAND2_X1 U1640 ( .A1(n1446), .A2(n917), .ZN(n1449) );
  FA_X1 U1641 ( .A(n1422), .B(n1421), .CI(n1420), .S(n1434) );
  NOR2_X1 U1642 ( .A1(n1449), .A2(n916), .ZN(n1423) );
  NOR2_X1 U1643 ( .A1(n1451), .A2(n1450), .ZN(n1452) );
  NOR2_X1 U1644 ( .A1(n915), .A2(n1452), .ZN(n1454) );
  NAND2_X1 U1645 ( .A1(n1423), .A2(n1454), .ZN(n1457) );
  NOR2_X1 U1646 ( .A1(n1424), .A2(n1457), .ZN(n1425) );
  NAND2_X1 U1647 ( .A1(n1602), .A2(n1425), .ZN(n1461) );
  NAND2_X1 U1648 ( .A1(n1427), .A2(n1426), .ZN(n1428) );
  OAI21_X1 U1649 ( .B1(n891), .B2(n1429), .A(n1428), .ZN(n1437) );
  NAND2_X1 U1650 ( .A1(n1432), .A2(n1431), .ZN(n1435) );
  OAI21_X1 U1651 ( .B1(n880), .B2(n1435), .A(n913), .ZN(n1436) );
  AOI21_X1 U1652 ( .B1(n1438), .B2(n1437), .A(n1436), .ZN(n1458) );
  XNOR2_X1 U1653 ( .A(n1442), .B(n1441), .ZN(n1447) );
  XNOR2_X1 U1654 ( .A(n1444), .B(n1443), .ZN(n1445) );
  AOI21_X1 U1655 ( .B1(n1447), .B2(n1446), .A(n1445), .ZN(n1448) );
  OAI21_X1 U1656 ( .B1(n914), .B2(n1449), .A(n1448), .ZN(n1455) );
  NOR2_X1 U1657 ( .A1(n912), .A2(n1452), .ZN(n1453) );
  AOI21_X1 U1658 ( .B1(n1455), .B2(n1454), .A(n1453), .ZN(n1456) );
  OAI21_X1 U1659 ( .B1(n1458), .B2(n1457), .A(n1456), .ZN(n1459) );
  INV_X1 U1660 ( .A(n1459), .ZN(n1460) );
  AND2_X2 U1661 ( .A1(n1461), .A2(n1460), .ZN(n1663) );
  AND2_X1 U1662 ( .A1(n1725), .A2(n1462), .ZN(n1463) );
  NAND2_X1 U1663 ( .A1(n1811), .A2(n1463), .ZN(n1592) );
  OAI211_X1 U1664 ( .C1(n1465), .C2(n1464), .A(n1663), .B(n1601), .ZN(n1466)
         );
  OAI21_X1 U1665 ( .B1(n1822), .B2(n1723), .A(n1466), .ZN(n596) );
  NOR3_X1 U1666 ( .A1(\ctrl_conv_output_inst/m_pre_valid_y ), .A2(n1836), .A3(
        n1467), .ZN(n1468) );
  NAND3_X1 U1667 ( .A1(\ctrl_conv_output_inst/cnt_conv [0]), .A2(
        \ctrl_conv_output_inst/cnt_conv [1]), .A3(n1468), .ZN(n1733) );
  NOR2_X1 U1668 ( .A1(n1837), .A2(n1733), .ZN(n1471) );
  INV_X1 U1669 ( .A(n1468), .ZN(n1730) );
  NAND2_X1 U1670 ( .A1(\ctrl_conv_output_inst/m_pre_pre_valid_y ), .A2(n1870), 
        .ZN(n1728) );
  OAI21_X1 U1671 ( .B1(n1841), .B2(n1728), .A(n1736), .ZN(n1731) );
  OAI21_X1 U1672 ( .B1(\ctrl_conv_output_inst/cnt_conv [1]), .B2(n1730), .A(
        n1731), .ZN(n1732) );
  AOI21_X1 U1673 ( .B1(n1468), .B2(n1837), .A(n1732), .ZN(n1469) );
  INV_X1 U1674 ( .A(n1469), .ZN(n1470) );
  MUX2_X1 U1675 ( .A(n1471), .B(n1470), .S(\ctrl_conv_output_inst/cnt_conv [3]), .Z(n878) );
  NAND2_X1 U1676 ( .A1(n1834), .A2(\fmem_inst/N12 ), .ZN(\fmem_inst/N13 ) );
  INV_X1 U1677 ( .A(n1476), .ZN(n1472) );
  NOR2_X2 U1678 ( .A1(n1473), .A2(n1472), .ZN(n1588) );
  OR2_X1 U1679 ( .A1(\mac_unit_inst/adder_reg [0]), .A2(
        \mac_unit_inst/x_mult_f_reg [0]), .ZN(n1474) );
  AND2_X1 U1680 ( .A1(n1474), .A2(n1482), .ZN(n1475) );
  NAND2_X1 U1681 ( .A1(n1588), .A2(n1475), .ZN(n1478) );
  OAI211_X1 U1682 ( .C1(n1591), .C2(n1868), .A(n1478), .B(n1589), .ZN(n595) );
  INV_X1 U1683 ( .A(n1479), .ZN(n1481) );
  NAND2_X1 U1684 ( .A1(n1481), .A2(n1480), .ZN(n1483) );
  XOR2_X1 U1685 ( .A(n1483), .B(n1482), .Z(n1484) );
  NAND2_X1 U1686 ( .A1(n1588), .A2(n1484), .ZN(n1485) );
  OAI211_X1 U1687 ( .C1(n1591), .C2(n1865), .A(n1485), .B(n1589), .ZN(n594) );
  INV_X1 U1688 ( .A(n1486), .ZN(n1493) );
  INV_X1 U1689 ( .A(n1492), .ZN(n1487) );
  NAND2_X1 U1690 ( .A1(n1487), .A2(n1491), .ZN(n1488) );
  XOR2_X1 U1691 ( .A(n1493), .B(n1488), .Z(n1489) );
  NAND2_X1 U1692 ( .A1(n1588), .A2(n1489), .ZN(n1490) );
  OAI211_X1 U1693 ( .C1(n1591), .C2(n1866), .A(n1490), .B(n1589), .ZN(n593) );
  OAI21_X1 U1694 ( .B1(n1493), .B2(n1492), .A(n1491), .ZN(n1498) );
  INV_X1 U1695 ( .A(n1494), .ZN(n1496) );
  NAND2_X1 U1696 ( .A1(n1496), .A2(n1495), .ZN(n1497) );
  XNOR2_X1 U1697 ( .A(n1498), .B(n1497), .ZN(n1499) );
  NAND2_X1 U1698 ( .A1(n1588), .A2(n1499), .ZN(n1500) );
  OAI211_X1 U1699 ( .C1(n1591), .C2(n1864), .A(n1500), .B(n1589), .ZN(n592) );
  INV_X1 U1700 ( .A(n1501), .ZN(n1518) );
  INV_X1 U1701 ( .A(n1502), .ZN(n1508) );
  NAND2_X1 U1702 ( .A1(n1508), .A2(n1506), .ZN(n1503) );
  XNOR2_X1 U1703 ( .A(n1518), .B(n1503), .ZN(n1504) );
  NAND2_X1 U1704 ( .A1(n1588), .A2(n1504), .ZN(n1505) );
  OAI211_X1 U1705 ( .C1(n1591), .C2(n1869), .A(n1505), .B(n1589), .ZN(n591) );
  INV_X1 U1706 ( .A(n1506), .ZN(n1507) );
  AOI21_X1 U1707 ( .B1(n1518), .B2(n1508), .A(n1507), .ZN(n1513) );
  INV_X1 U1708 ( .A(n1509), .ZN(n1511) );
  NAND2_X1 U1709 ( .A1(n1511), .A2(n1510), .ZN(n1512) );
  XOR2_X1 U1710 ( .A(n1513), .B(n1512), .Z(n1514) );
  NAND2_X1 U1711 ( .A1(n1588), .A2(n1514), .ZN(n1515) );
  OAI211_X1 U1712 ( .C1(n1591), .C2(n1871), .A(n1515), .B(n1589), .ZN(n590) );
  AOI21_X1 U1713 ( .B1(n1518), .B2(n1517), .A(n1516), .ZN(n1525) );
  INV_X1 U1714 ( .A(n1524), .ZN(n1519) );
  NAND2_X1 U1715 ( .A1(n1519), .A2(n1523), .ZN(n1520) );
  XOR2_X1 U1716 ( .A(n1525), .B(n1520), .Z(n1521) );
  NAND2_X1 U1717 ( .A1(n1588), .A2(n1521), .ZN(n1522) );
  OAI211_X1 U1718 ( .C1(n1591), .C2(n1867), .A(n1522), .B(n1589), .ZN(n589) );
  OAI21_X1 U1719 ( .B1(n1525), .B2(n1524), .A(n1523), .ZN(n1530) );
  INV_X1 U1720 ( .A(n1526), .ZN(n1528) );
  NAND2_X1 U1721 ( .A1(n1528), .A2(n1527), .ZN(n1529) );
  XNOR2_X1 U1722 ( .A(n1530), .B(n1529), .ZN(n1531) );
  NAND2_X1 U1723 ( .A1(n1588), .A2(n1531), .ZN(n1532) );
  OAI211_X1 U1724 ( .C1(n1591), .C2(n1872), .A(n1532), .B(n1589), .ZN(n588) );
  INV_X1 U1725 ( .A(n1533), .ZN(n1586) );
  OAI21_X1 U1726 ( .B1(n1586), .B2(n1582), .A(n1583), .ZN(n1538) );
  INV_X1 U1727 ( .A(n1534), .ZN(n1536) );
  NAND2_X1 U1728 ( .A1(n1536), .A2(n1535), .ZN(n1537) );
  XNOR2_X1 U1729 ( .A(n1538), .B(n1537), .ZN(n1539) );
  NAND2_X1 U1730 ( .A1(n1588), .A2(n1539), .ZN(n1540) );
  OAI211_X1 U1731 ( .C1(n1591), .C2(n1844), .A(n1540), .B(n1589), .ZN(n586) );
  INV_X1 U1732 ( .A(n1541), .ZN(n1544) );
  INV_X1 U1733 ( .A(n1542), .ZN(n1543) );
  OAI21_X1 U1734 ( .B1(n1586), .B2(n1544), .A(n1543), .ZN(n1552) );
  INV_X1 U1735 ( .A(n1545), .ZN(n1551) );
  NAND2_X1 U1736 ( .A1(n1551), .A2(n1549), .ZN(n1546) );
  XNOR2_X1 U1737 ( .A(n1552), .B(n1546), .ZN(n1547) );
  NAND2_X1 U1738 ( .A1(n1588), .A2(n1547), .ZN(n1548) );
  OAI211_X1 U1739 ( .C1(n1591), .C2(n1845), .A(n1548), .B(n1589), .ZN(n585) );
  INV_X1 U1740 ( .A(n1549), .ZN(n1550) );
  AOI21_X1 U1741 ( .B1(n1552), .B2(n1551), .A(n1550), .ZN(n1557) );
  INV_X1 U1742 ( .A(n1553), .ZN(n1555) );
  NAND2_X1 U1743 ( .A1(n1555), .A2(n1554), .ZN(n1556) );
  XOR2_X1 U1744 ( .A(n1557), .B(n1556), .Z(n1558) );
  NAND2_X1 U1745 ( .A1(n1588), .A2(n1558), .ZN(n1559) );
  OAI211_X1 U1746 ( .C1(n1591), .C2(n1873), .A(n1559), .B(n1589), .ZN(n584) );
  INV_X1 U1747 ( .A(n1568), .ZN(n1562) );
  INV_X1 U1748 ( .A(n1560), .ZN(n1567) );
  NAND2_X1 U1749 ( .A1(n1567), .A2(n1565), .ZN(n1561) );
  XOR2_X1 U1750 ( .A(n1562), .B(n1561), .Z(n1563) );
  NAND2_X1 U1751 ( .A1(n1588), .A2(n1563), .ZN(n1564) );
  OAI211_X1 U1752 ( .C1(n1591), .C2(n1846), .A(n1564), .B(n1589), .ZN(n583) );
  INV_X1 U1753 ( .A(n1565), .ZN(n1566) );
  AOI21_X1 U1754 ( .B1(n1568), .B2(n1567), .A(n1566), .ZN(n1573) );
  INV_X1 U1755 ( .A(n1569), .ZN(n1571) );
  NAND2_X1 U1756 ( .A1(n1571), .A2(n1570), .ZN(n1572) );
  XOR2_X1 U1757 ( .A(n1573), .B(n1572), .Z(n1574) );
  NAND2_X1 U1758 ( .A1(n1588), .A2(n1574), .ZN(n1575) );
  OAI211_X1 U1759 ( .C1(n1591), .C2(n1874), .A(n1575), .B(n1589), .ZN(n582) );
  NAND2_X1 U1760 ( .A1(n1577), .A2(n1576), .ZN(n1578) );
  XNOR2_X1 U1761 ( .A(n1579), .B(n1578), .ZN(n1580) );
  NAND2_X1 U1762 ( .A1(n1588), .A2(n1580), .ZN(n1581) );
  OAI211_X1 U1763 ( .C1(n1591), .C2(n1847), .A(n1581), .B(n1589), .ZN(n581) );
  INV_X1 U1764 ( .A(n1582), .ZN(n1584) );
  NAND2_X1 U1765 ( .A1(n1584), .A2(n1583), .ZN(n1585) );
  XOR2_X1 U1766 ( .A(n1586), .B(n1585), .Z(n1587) );
  NAND2_X1 U1767 ( .A1(n1588), .A2(n1587), .ZN(n1590) );
  OAI211_X1 U1768 ( .C1(n1591), .C2(n1843), .A(n1590), .B(n1589), .ZN(n587) );
  INV_X1 U1769 ( .A(n1592), .ZN(n1601) );
  NAND2_X1 U1770 ( .A1(n1593), .A2(n1601), .ZN(n1604) );
  NOR2_X1 U1771 ( .A1(n1594), .A2(n1595), .ZN(n1596) );
  NAND2_X1 U1772 ( .A1(n1597), .A2(n1596), .ZN(n1599) );
  NOR2_X1 U1773 ( .A1(n1599), .A2(n1598), .ZN(n1600) );
  NAND3_X1 U1774 ( .A1(n1602), .A2(n1601), .A3(n1600), .ZN(n1603) );
  NAND2_X1 U1775 ( .A1(n1603), .A2(n1604), .ZN(n1620) );
  BUF_X1 U1776 ( .A(n1620), .Z(n1704) );
  NOR2_X1 U1777 ( .A1(n1605), .A2(n1824), .ZN(n1606) );
  NAND2_X1 U1778 ( .A1(n1704), .A2(n1606), .ZN(n1607) );
  OR2_X2 U1779 ( .A1(n1663), .A2(n1592), .ZN(n1721) );
  OAI211_X1 U1780 ( .C1(n1723), .C2(n2118), .A(n1607), .B(n1721), .ZN(n611) );
  BUF_X1 U1781 ( .A(n902), .Z(n1679) );
  OR2_X1 U1782 ( .A1(n1608), .A2(n884), .ZN(n1609) );
  AND2_X1 U1783 ( .A1(n1609), .A2(n1616), .ZN(n1610) );
  NAND2_X1 U1784 ( .A1(n905), .A2(n1610), .ZN(n1611) );
  OR2_X2 U1785 ( .A1(n1663), .A2(n1592), .ZN(n1705) );
  OAI211_X1 U1786 ( .C1(n1723), .C2(n2119), .A(n1611), .B(n1705), .ZN(n610) );
  OR2_X1 U1787 ( .A1(n1613), .A2(n1612), .ZN(n1615) );
  NAND2_X1 U1788 ( .A1(n1615), .A2(n1614), .ZN(n1617) );
  XOR2_X1 U1789 ( .A(n1617), .B(n1616), .Z(n1618) );
  NAND2_X1 U1790 ( .A1(n1679), .A2(n1618), .ZN(n1619) );
  OAI211_X1 U1791 ( .C1(n1723), .C2(n2120), .A(n1619), .B(n1721), .ZN(n609) );
  BUF_X1 U1792 ( .A(n902), .Z(n1720) );
  NAND2_X1 U1793 ( .A1(n1622), .A2(n1621), .ZN(n1623) );
  XNOR2_X1 U1794 ( .A(n1624), .B(n1623), .ZN(n1625) );
  NAND2_X1 U1795 ( .A1(n904), .A2(n1625), .ZN(n1626) );
  OAI211_X1 U1796 ( .C1(n1723), .C2(n2121), .A(n1626), .B(n1705), .ZN(n608) );
  INV_X1 U1797 ( .A(n1627), .ZN(n1629) );
  NAND2_X1 U1798 ( .A1(n1629), .A2(n1628), .ZN(n1631) );
  XOR2_X1 U1799 ( .A(n1631), .B(n1630), .Z(n1632) );
  NAND2_X1 U1800 ( .A1(n1720), .A2(n1632), .ZN(n1633) );
  OAI211_X1 U1801 ( .C1(n1723), .C2(n2122), .A(n1633), .B(n1721), .ZN(n607) );
  XNOR2_X1 U1802 ( .A(n1638), .B(n885), .ZN(n1639) );
  NAND2_X1 U1803 ( .A1(n1720), .A2(n1639), .ZN(n1640) );
  OAI211_X1 U1804 ( .C1(n1723), .C2(n2123), .A(n1640), .B(n1705), .ZN(n606) );
  INV_X1 U1805 ( .A(n893), .ZN(n1644) );
  NAND2_X1 U1806 ( .A1(n1644), .A2(n1643), .ZN(n1645) );
  XOR2_X1 U1807 ( .A(n1641), .B(n1645), .Z(n1646) );
  NAND2_X1 U1808 ( .A1(n905), .A2(n1646), .ZN(n1647) );
  OAI211_X1 U1809 ( .C1(n1723), .C2(n2124), .A(n1647), .B(n1721), .ZN(n605) );
  INV_X1 U1810 ( .A(n1648), .ZN(n1650) );
  NAND2_X1 U1811 ( .A1(n1650), .A2(n1649), .ZN(n1653) );
  XNOR2_X1 U1812 ( .A(n1653), .B(n1652), .ZN(n1654) );
  NAND2_X1 U1813 ( .A1(n905), .A2(n1654), .ZN(n1655) );
  OAI211_X1 U1814 ( .C1(n1723), .C2(n2125), .A(n1655), .B(n1705), .ZN(n604) );
  INV_X1 U1815 ( .A(n1657), .ZN(n1659) );
  NAND2_X1 U1816 ( .A1(n1659), .A2(n1658), .ZN(n1660) );
  XOR2_X1 U1817 ( .A(n1661), .B(n1660), .Z(n1662) );
  NAND2_X1 U1818 ( .A1(n1704), .A2(n1662), .ZN(n1664) );
  OR2_X2 U1819 ( .A1(n1663), .A2(n1592), .ZN(n1695) );
  OAI211_X1 U1820 ( .C1(n1723), .C2(n2126), .A(n1664), .B(n1695), .ZN(n603) );
  INV_X1 U1821 ( .A(n1671), .ZN(n1665) );
  NAND2_X1 U1822 ( .A1(n1665), .A2(n883), .ZN(n1667) );
  INV_X1 U1823 ( .A(n1666), .ZN(n1672) );
  XOR2_X1 U1824 ( .A(n1667), .B(n1672), .Z(n1668) );
  NAND2_X1 U1825 ( .A1(n904), .A2(n1668), .ZN(n1669) );
  OAI211_X1 U1826 ( .C1(n1723), .C2(n2127), .A(n1669), .B(n1695), .ZN(n602) );
  OAI21_X1 U1827 ( .B1(n1672), .B2(n1671), .A(n883), .ZN(n1677) );
  INV_X1 U1828 ( .A(n1673), .ZN(n1675) );
  NAND2_X1 U1829 ( .A1(n1675), .A2(n1674), .ZN(n1676) );
  XNOR2_X1 U1830 ( .A(n1677), .B(n1676), .ZN(n1678) );
  NAND2_X1 U1831 ( .A1(n1720), .A2(n1678), .ZN(n1680) );
  OAI211_X1 U1832 ( .C1(n1723), .C2(n2128), .A(n1680), .B(n1695), .ZN(n601) );
  INV_X1 U1833 ( .A(n1681), .ZN(n1712) );
  INV_X1 U1834 ( .A(n1682), .ZN(n1688) );
  INV_X1 U1835 ( .A(n1683), .ZN(n1687) );
  NAND2_X1 U1836 ( .A1(n1688), .A2(n1683), .ZN(n1684) );
  XNOR2_X1 U1837 ( .A(n1712), .B(n1684), .ZN(n1685) );
  NAND2_X1 U1838 ( .A1(n1679), .A2(n1685), .ZN(n1686) );
  OAI211_X1 U1839 ( .C1(n1723), .C2(n2129), .A(n1686), .B(n1695), .ZN(n600) );
  AOI21_X1 U1840 ( .B1(n1712), .B2(n1688), .A(n1687), .ZN(n1693) );
  INV_X1 U1841 ( .A(n898), .ZN(n1691) );
  NAND2_X1 U1842 ( .A1(n1691), .A2(n1690), .ZN(n1692) );
  XOR2_X1 U1843 ( .A(n1693), .B(n1692), .Z(n1694) );
  NAND2_X1 U1844 ( .A1(n904), .A2(n1694), .ZN(n1696) );
  OAI211_X1 U1845 ( .C1(n1723), .C2(n2130), .A(n1696), .B(n1695), .ZN(n599) );
  INV_X1 U1846 ( .A(n900), .ZN(n1708) );
  INV_X1 U1847 ( .A(n1698), .ZN(n1710) );
  INV_X1 U1848 ( .A(n1710), .ZN(n1699) );
  AOI21_X1 U1849 ( .B1(n1712), .B2(n900), .A(n1699), .ZN(n1702) );
  INV_X1 U1850 ( .A(n1700), .ZN(n1707) );
  NAND2_X1 U1851 ( .A1(n1707), .A2(n1709), .ZN(n1701) );
  XOR2_X1 U1852 ( .A(n1702), .B(n1701), .Z(n1703) );
  NAND2_X1 U1853 ( .A1(n1679), .A2(n1703), .ZN(n1706) );
  OAI211_X1 U1854 ( .C1(n1723), .C2(n2131), .A(n1706), .B(n1705), .ZN(n598) );
  NOR2_X1 U1855 ( .A1(n1708), .A2(n901), .ZN(n1713) );
  OAI21_X1 U1856 ( .B1(n1710), .B2(n901), .A(n1709), .ZN(n1711) );
  AOI21_X1 U1857 ( .B1(n1713), .B2(n1712), .A(n1711), .ZN(n1718) );
  INV_X1 U1858 ( .A(n1714), .ZN(n1716) );
  NAND2_X1 U1859 ( .A1(n1716), .A2(n1715), .ZN(n1717) );
  XOR2_X1 U1860 ( .A(n1718), .B(n1717), .Z(n1719) );
  NAND2_X1 U1861 ( .A1(n1704), .A2(n1719), .ZN(n1722) );
  OAI211_X1 U1862 ( .C1(n1723), .C2(n2132), .A(n1722), .B(n1721), .ZN(n597) );
  NAND2_X1 U1864 ( .A1(\ctrl_conv_output_inst/cnt_conv [0]), .A2(n1840), .ZN(
        n1729) );
  NAND4_X1 U1865 ( .A1(n1727), .A2(\ctrl_conv_output_inst/cnt_conv [2]), .A3(
        \ctrl_conv_output_inst/cnt_conv [3]), .A4(n1812), .ZN(n1724) );
  NOR2_X1 U1866 ( .A1(n1729), .A2(n1724), .ZN(\ctrl_conv_output_inst/N74 ) );
  NOR2_X1 U1867 ( .A1(reset), .A2(s_ready_x), .ZN(N19) );
  NAND3_X1 U1868 ( .A1(n1725), .A2(\fmem_inst/N12 ), .A3(\fmem_inst/N14 ), 
        .ZN(n1726) );
  AOI221_X1 U1869 ( .B1(n1727), .B2(\ctrl_conv_output_inst/m_pre_pre_valid_y ), 
        .C1(n1726), .C2(n1836), .A(reset), .ZN(n879) );
  AOI21_X1 U1870 ( .B1(n1841), .B2(n1728), .A(n1731), .ZN(n877) );
  OAI22_X1 U1871 ( .A1(n1840), .A2(n1731), .B1(n1730), .B2(n1729), .ZN(n876)
         );
  INV_X1 U1872 ( .A(n1732), .ZN(n1734) );
  AOI22_X1 U1873 ( .A1(\ctrl_conv_output_inst/cnt_conv [2]), .A2(n1734), .B1(
        n1733), .B2(n1837), .ZN(n875) );
  OAI21_X1 U1874 ( .B1(n1810), .B2(n2116), .A(n1736), .ZN(n873) );
  NAND2_X1 U1875 ( .A1(n1743), .A2(\ctrl_conv_output_inst/cnt_conv [0]), .ZN(
        n1737) );
  OAI221_X1 U1876 ( .B1(xmem_addr[0]), .B2(n1745), .C1(n1833), .C2(n1738), .A(
        n1737), .ZN(n872) );
  AOI22_X1 U1877 ( .A1(xmem_addr[1]), .A2(n1739), .B1(n1743), .B2(
        \ctrl_conv_output_inst/cnt_conv [1]), .ZN(n1740) );
  OAI221_X1 U1878 ( .B1(n1745), .B2(n1752), .C1(n1745), .C2(n1741), .A(n1740), 
        .ZN(n871) );
  AOI22_X1 U1879 ( .A1(\ctrl_conv_output_inst/cnt_conv [3]), .A2(n1743), .B1(
        xmem_addr[3]), .B2(n1742), .ZN(n1744) );
  OAI221_X1 U1880 ( .B1(n1745), .B2(n1776), .C1(n1745), .C2(n1767), .A(n1744), 
        .ZN(n869) );
  NOR2_X2 U1881 ( .A1(n1753), .A2(n1782), .ZN(n1748) );
  INV_X1 U1882 ( .A(s_data_in_x[0]), .ZN(n1793) );
  AOI22_X1 U1883 ( .A1(n1748), .A2(n1793), .B1(n2036), .B2(n1747), .ZN(n868)
         );
  INV_X1 U1884 ( .A(s_data_in_x[1]), .ZN(n1794) );
  AOI22_X1 U1885 ( .A1(n1748), .A2(n1794), .B1(n2037), .B2(n1747), .ZN(n867)
         );
  INV_X1 U1886 ( .A(s_data_in_x[2]), .ZN(n1795) );
  AOI22_X1 U1887 ( .A1(n1748), .A2(n1795), .B1(n2038), .B2(n1747), .ZN(n866)
         );
  INV_X1 U1888 ( .A(s_data_in_x[3]), .ZN(n1796) );
  AOI22_X1 U1889 ( .A1(n1748), .A2(n1796), .B1(n2039), .B2(n1747), .ZN(n865)
         );
  INV_X1 U1890 ( .A(s_data_in_x[4]), .ZN(n1797) );
  AOI22_X1 U1891 ( .A1(n1748), .A2(n1797), .B1(n2040), .B2(n1747), .ZN(n864)
         );
  INV_X1 U1892 ( .A(s_data_in_x[5]), .ZN(n1798) );
  AOI22_X1 U1893 ( .A1(n1748), .A2(n1798), .B1(n2041), .B2(n1747), .ZN(n863)
         );
  INV_X1 U1894 ( .A(s_data_in_x[6]), .ZN(n1799) );
  AOI22_X1 U1895 ( .A1(n1748), .A2(n1799), .B1(n2042), .B2(n1747), .ZN(n862)
         );
  INV_X1 U1896 ( .A(s_data_in_x[7]), .ZN(n1800) );
  AOI22_X1 U1897 ( .A1(n1748), .A2(n1800), .B1(n2043), .B2(n1747), .ZN(n861)
         );
  INV_X1 U1898 ( .A(s_data_in_x[8]), .ZN(n1801) );
  AOI22_X1 U1899 ( .A1(n1748), .A2(n1801), .B1(n2044), .B2(n1747), .ZN(n860)
         );
  INV_X1 U1900 ( .A(s_data_in_x[9]), .ZN(n1802) );
  AOI22_X1 U1901 ( .A1(n1748), .A2(n1802), .B1(n2045), .B2(n1747), .ZN(n859)
         );
  INV_X1 U1902 ( .A(s_data_in_x[10]), .ZN(n1803) );
  AOI22_X1 U1903 ( .A1(n1748), .A2(n1803), .B1(n2046), .B2(n1747), .ZN(n858)
         );
  INV_X1 U1904 ( .A(s_data_in_x[11]), .ZN(n1804) );
  AOI22_X1 U1905 ( .A1(n1748), .A2(n1804), .B1(n2047), .B2(n1747), .ZN(n857)
         );
  INV_X1 U1906 ( .A(s_data_in_x[12]), .ZN(n1805) );
  AOI22_X1 U1907 ( .A1(n1748), .A2(n1805), .B1(n2048), .B2(n1747), .ZN(n856)
         );
  INV_X1 U1908 ( .A(s_data_in_x[13]), .ZN(n1806) );
  AOI22_X1 U1909 ( .A1(n1748), .A2(n1806), .B1(n2049), .B2(n1747), .ZN(n855)
         );
  INV_X1 U1910 ( .A(s_data_in_x[14]), .ZN(n1807) );
  AOI22_X1 U1911 ( .A1(n1748), .A2(n1807), .B1(n2050), .B2(n1747), .ZN(n854)
         );
  INV_X1 U1912 ( .A(s_data_in_x[15]), .ZN(n1809) );
  AOI22_X1 U1913 ( .A1(n1748), .A2(n1809), .B1(n2051), .B2(n1747), .ZN(n853)
         );
  AOI22_X1 U1914 ( .A1(n1751), .A2(n1793), .B1(n1955), .B2(n1750), .ZN(n852)
         );
  AOI22_X1 U1915 ( .A1(n1751), .A2(n1794), .B1(n1956), .B2(n1750), .ZN(n851)
         );
  AOI22_X1 U1916 ( .A1(n1751), .A2(n1795), .B1(n1957), .B2(n1750), .ZN(n850)
         );
  AOI22_X1 U1917 ( .A1(n1751), .A2(n1796), .B1(n1958), .B2(n1750), .ZN(n849)
         );
  AOI22_X1 U1918 ( .A1(n1751), .A2(n1797), .B1(n1959), .B2(n1750), .ZN(n848)
         );
  AOI22_X1 U1919 ( .A1(n1751), .A2(n1798), .B1(n1960), .B2(n1750), .ZN(n847)
         );
  AOI22_X1 U1920 ( .A1(n1751), .A2(n1799), .B1(n1961), .B2(n1750), .ZN(n846)
         );
  AOI22_X1 U1921 ( .A1(n1751), .A2(n1800), .B1(n1962), .B2(n1750), .ZN(n845)
         );
  AOI22_X1 U1922 ( .A1(n1751), .A2(n1801), .B1(n1963), .B2(n1750), .ZN(n844)
         );
  AOI22_X1 U1923 ( .A1(n1751), .A2(n1802), .B1(n1964), .B2(n1750), .ZN(n843)
         );
  AOI22_X1 U1924 ( .A1(n1751), .A2(n1803), .B1(n1965), .B2(n1750), .ZN(n842)
         );
  AOI22_X1 U1925 ( .A1(n1751), .A2(n1804), .B1(n1966), .B2(n1750), .ZN(n841)
         );
  AOI22_X1 U1926 ( .A1(n1751), .A2(n1805), .B1(n1967), .B2(n1750), .ZN(n840)
         );
  AOI22_X1 U1927 ( .A1(n1751), .A2(n1806), .B1(n1968), .B2(n1750), .ZN(n839)
         );
  AOI22_X1 U1928 ( .A1(n1751), .A2(n1807), .B1(n1969), .B2(n1750), .ZN(n838)
         );
  AOI22_X1 U1929 ( .A1(n1751), .A2(n1809), .B1(n1970), .B2(n1750), .ZN(n837)
         );
  NOR2_X2 U1930 ( .A1(n1753), .A2(n1789), .ZN(n1755) );
  AOI22_X1 U1931 ( .A1(n1755), .A2(n1793), .B1(n2052), .B2(n1754), .ZN(n836)
         );
  AOI22_X1 U1932 ( .A1(n1755), .A2(n1794), .B1(n2053), .B2(n1754), .ZN(n835)
         );
  AOI22_X1 U1933 ( .A1(n1755), .A2(n1795), .B1(n2054), .B2(n1754), .ZN(n834)
         );
  AOI22_X1 U1934 ( .A1(n1755), .A2(n1796), .B1(n2055), .B2(n1754), .ZN(n833)
         );
  AOI22_X1 U1935 ( .A1(n1755), .A2(n1797), .B1(n2056), .B2(n1754), .ZN(n832)
         );
  AOI22_X1 U1936 ( .A1(n1755), .A2(n1798), .B1(n2057), .B2(n1754), .ZN(n831)
         );
  AOI22_X1 U1937 ( .A1(n1755), .A2(n1799), .B1(n2058), .B2(n1754), .ZN(n830)
         );
  AOI22_X1 U1938 ( .A1(n1755), .A2(n1800), .B1(n2059), .B2(n1754), .ZN(n829)
         );
  AOI22_X1 U1939 ( .A1(n1755), .A2(n1801), .B1(n2060), .B2(n1754), .ZN(n828)
         );
  AOI22_X1 U1940 ( .A1(n1755), .A2(n1802), .B1(n2061), .B2(n1754), .ZN(n827)
         );
  AOI22_X1 U1941 ( .A1(n1755), .A2(n1803), .B1(n2062), .B2(n1754), .ZN(n826)
         );
  AOI22_X1 U1942 ( .A1(n1755), .A2(n1804), .B1(n2063), .B2(n1754), .ZN(n825)
         );
  AOI22_X1 U1943 ( .A1(n1755), .A2(n1805), .B1(n2064), .B2(n1754), .ZN(n824)
         );
  AOI22_X1 U1944 ( .A1(n1755), .A2(n1806), .B1(n2065), .B2(n1754), .ZN(n823)
         );
  AOI22_X1 U1945 ( .A1(n1755), .A2(n1807), .B1(n2066), .B2(n1754), .ZN(n822)
         );
  AOI22_X1 U1946 ( .A1(n1755), .A2(n1809), .B1(n2067), .B2(n1754), .ZN(n821)
         );
  AOI22_X1 U1947 ( .A1(n1758), .A2(n1793), .B1(n1971), .B2(n1757), .ZN(n820)
         );
  AOI22_X1 U1948 ( .A1(n1758), .A2(n1794), .B1(n1972), .B2(n1757), .ZN(n819)
         );
  AOI22_X1 U1949 ( .A1(n1758), .A2(n1795), .B1(n1973), .B2(n1757), .ZN(n818)
         );
  AOI22_X1 U1950 ( .A1(n1758), .A2(n1796), .B1(n1974), .B2(n1757), .ZN(n817)
         );
  AOI22_X1 U1951 ( .A1(n1758), .A2(n1797), .B1(n1975), .B2(n1757), .ZN(n816)
         );
  AOI22_X1 U1952 ( .A1(n1758), .A2(n1798), .B1(n1976), .B2(n1757), .ZN(n815)
         );
  AOI22_X1 U1953 ( .A1(n1758), .A2(n1799), .B1(n1977), .B2(n1757), .ZN(n814)
         );
  AOI22_X1 U1954 ( .A1(n1758), .A2(n1800), .B1(n1978), .B2(n1757), .ZN(n813)
         );
  AOI22_X1 U1955 ( .A1(n1758), .A2(n1801), .B1(n1979), .B2(n1757), .ZN(n812)
         );
  AOI22_X1 U1956 ( .A1(n1758), .A2(n1802), .B1(n1980), .B2(n1757), .ZN(n811)
         );
  AOI22_X1 U1957 ( .A1(n1758), .A2(n1803), .B1(n1981), .B2(n1757), .ZN(n810)
         );
  AOI22_X1 U1958 ( .A1(n1758), .A2(n1804), .B1(n1982), .B2(n1757), .ZN(n809)
         );
  AOI22_X1 U1959 ( .A1(n1758), .A2(n1805), .B1(n1983), .B2(n1757), .ZN(n808)
         );
  AOI22_X1 U1960 ( .A1(n1758), .A2(n1806), .B1(n1984), .B2(n1757), .ZN(n807)
         );
  AOI22_X1 U1961 ( .A1(n1758), .A2(n1807), .B1(n1985), .B2(n1757), .ZN(n806)
         );
  AOI22_X1 U1962 ( .A1(n1758), .A2(n1809), .B1(n1986), .B2(n1757), .ZN(n805)
         );
  NOR2_X2 U1963 ( .A1(n1764), .A2(n1782), .ZN(n1760) );
  AOI22_X1 U1964 ( .A1(n1760), .A2(n1793), .B1(n2068), .B2(n1759), .ZN(n804)
         );
  AOI22_X1 U1965 ( .A1(n1760), .A2(n1794), .B1(n2069), .B2(n1759), .ZN(n803)
         );
  AOI22_X1 U1966 ( .A1(n1760), .A2(n1795), .B1(n2070), .B2(n1759), .ZN(n802)
         );
  AOI22_X1 U1967 ( .A1(n1760), .A2(n1796), .B1(n2071), .B2(n1759), .ZN(n801)
         );
  AOI22_X1 U1968 ( .A1(n1760), .A2(n1797), .B1(n2072), .B2(n1759), .ZN(n800)
         );
  AOI22_X1 U1969 ( .A1(n1760), .A2(n1798), .B1(n2073), .B2(n1759), .ZN(n799)
         );
  AOI22_X1 U1970 ( .A1(n1760), .A2(n1799), .B1(n2074), .B2(n1759), .ZN(n798)
         );
  AOI22_X1 U1971 ( .A1(n1760), .A2(n1800), .B1(n2075), .B2(n1759), .ZN(n797)
         );
  AOI22_X1 U1972 ( .A1(n1760), .A2(n1801), .B1(n2076), .B2(n1759), .ZN(n796)
         );
  AOI22_X1 U1973 ( .A1(n1760), .A2(n1802), .B1(n2077), .B2(n1759), .ZN(n795)
         );
  AOI22_X1 U1974 ( .A1(n1760), .A2(n1803), .B1(n2078), .B2(n1759), .ZN(n794)
         );
  AOI22_X1 U1975 ( .A1(n1760), .A2(n1804), .B1(n2079), .B2(n1759), .ZN(n793)
         );
  AOI22_X1 U1976 ( .A1(n1760), .A2(n1805), .B1(n2080), .B2(n1759), .ZN(n792)
         );
  AOI22_X1 U1977 ( .A1(n1760), .A2(n1806), .B1(n2081), .B2(n1759), .ZN(n791)
         );
  AOI22_X1 U1978 ( .A1(n1760), .A2(n1807), .B1(n2082), .B2(n1759), .ZN(n790)
         );
  AOI22_X1 U1979 ( .A1(n1760), .A2(n1809), .B1(n2083), .B2(n1759), .ZN(n789)
         );
  AOI22_X1 U1980 ( .A1(n1763), .A2(n1793), .B1(n1987), .B2(n1762), .ZN(n788)
         );
  AOI22_X1 U1981 ( .A1(n1763), .A2(n1794), .B1(n1988), .B2(n1762), .ZN(n787)
         );
  AOI22_X1 U1982 ( .A1(n1763), .A2(n1795), .B1(n1989), .B2(n1762), .ZN(n786)
         );
  AOI22_X1 U1983 ( .A1(n1763), .A2(n1796), .B1(n1990), .B2(n1762), .ZN(n785)
         );
  AOI22_X1 U1984 ( .A1(n1763), .A2(n1797), .B1(n1991), .B2(n1762), .ZN(n784)
         );
  AOI22_X1 U1985 ( .A1(n1763), .A2(n1798), .B1(n1992), .B2(n1762), .ZN(n783)
         );
  AOI22_X1 U1986 ( .A1(n1763), .A2(n1799), .B1(n1993), .B2(n1762), .ZN(n782)
         );
  AOI22_X1 U1987 ( .A1(n1763), .A2(n1800), .B1(n1994), .B2(n1762), .ZN(n781)
         );
  AOI22_X1 U1988 ( .A1(n1763), .A2(n1801), .B1(n1995), .B2(n1762), .ZN(n780)
         );
  AOI22_X1 U1989 ( .A1(n1763), .A2(n1802), .B1(n1996), .B2(n1762), .ZN(n779)
         );
  AOI22_X1 U1990 ( .A1(n1763), .A2(n1803), .B1(n1997), .B2(n1762), .ZN(n778)
         );
  AOI22_X1 U1991 ( .A1(n1763), .A2(n1804), .B1(n1998), .B2(n1762), .ZN(n777)
         );
  AOI22_X1 U1992 ( .A1(n1763), .A2(n1805), .B1(n1999), .B2(n1762), .ZN(n776)
         );
  AOI22_X1 U1993 ( .A1(n1763), .A2(n1806), .B1(n2000), .B2(n1762), .ZN(n775)
         );
  AOI22_X1 U1994 ( .A1(n1763), .A2(n1807), .B1(n2001), .B2(n1762), .ZN(n774)
         );
  AOI22_X1 U1995 ( .A1(n1763), .A2(n1809), .B1(n2002), .B2(n1762), .ZN(n773)
         );
  NOR2_X2 U1996 ( .A1(n1764), .A2(n1789), .ZN(n1766) );
  AOI22_X1 U1997 ( .A1(n1766), .A2(n1793), .B1(n1939), .B2(n1765), .ZN(n772)
         );
  AOI22_X1 U1998 ( .A1(n1766), .A2(n1794), .B1(n1940), .B2(n1765), .ZN(n771)
         );
  AOI22_X1 U1999 ( .A1(n1766), .A2(n1795), .B1(n1941), .B2(n1765), .ZN(n770)
         );
  AOI22_X1 U2000 ( .A1(n1766), .A2(n1796), .B1(n1942), .B2(n1765), .ZN(n769)
         );
  AOI22_X1 U2001 ( .A1(n1766), .A2(n1797), .B1(n1943), .B2(n1765), .ZN(n768)
         );
  AOI22_X1 U2002 ( .A1(n1766), .A2(n1798), .B1(n1944), .B2(n1765), .ZN(n767)
         );
  AOI22_X1 U2003 ( .A1(n1766), .A2(n1799), .B1(n1945), .B2(n1765), .ZN(n766)
         );
  AOI22_X1 U2004 ( .A1(n1766), .A2(n1800), .B1(n1946), .B2(n1765), .ZN(n765)
         );
  AOI22_X1 U2005 ( .A1(n1766), .A2(n1801), .B1(n1947), .B2(n1765), .ZN(n764)
         );
  AOI22_X1 U2006 ( .A1(n1766), .A2(n1802), .B1(n1948), .B2(n1765), .ZN(n763)
         );
  AOI22_X1 U2007 ( .A1(n1766), .A2(n1803), .B1(n1949), .B2(n1765), .ZN(n762)
         );
  AOI22_X1 U2008 ( .A1(n1766), .A2(n1804), .B1(n1950), .B2(n1765), .ZN(n761)
         );
  AOI22_X1 U2009 ( .A1(n1766), .A2(n1805), .B1(n1951), .B2(n1765), .ZN(n760)
         );
  AOI22_X1 U2010 ( .A1(n1766), .A2(n1806), .B1(n1952), .B2(n1765), .ZN(n759)
         );
  AOI22_X1 U2011 ( .A1(n1766), .A2(n1807), .B1(n1953), .B2(n1765), .ZN(n758)
         );
  AOI22_X1 U2012 ( .A1(n1766), .A2(n1809), .B1(n1954), .B2(n1765), .ZN(n757)
         );
  NOR2_X2 U2013 ( .A1(n1768), .A2(n1767), .ZN(n1770) );
  AOI22_X1 U2014 ( .A1(n1770), .A2(n1793), .B1(n1848), .B2(n1769), .ZN(n756)
         );
  AOI22_X1 U2015 ( .A1(n1770), .A2(n1794), .B1(n1849), .B2(n1769), .ZN(n755)
         );
  AOI22_X1 U2016 ( .A1(n1770), .A2(n1795), .B1(n1850), .B2(n1769), .ZN(n754)
         );
  AOI22_X1 U2017 ( .A1(n1770), .A2(n1796), .B1(n1851), .B2(n1769), .ZN(n753)
         );
  AOI22_X1 U2018 ( .A1(n1770), .A2(n1797), .B1(n1852), .B2(n1769), .ZN(n752)
         );
  AOI22_X1 U2019 ( .A1(n1770), .A2(n1798), .B1(n1853), .B2(n1769), .ZN(n751)
         );
  AOI22_X1 U2020 ( .A1(n1770), .A2(n1799), .B1(n1854), .B2(n1769), .ZN(n750)
         );
  AOI22_X1 U2021 ( .A1(n1770), .A2(n1800), .B1(n1855), .B2(n1769), .ZN(n749)
         );
  AOI22_X1 U2022 ( .A1(n1770), .A2(n1801), .B1(n1856), .B2(n1769), .ZN(n748)
         );
  AOI22_X1 U2023 ( .A1(n1770), .A2(n1802), .B1(n1857), .B2(n1769), .ZN(n747)
         );
  AOI22_X1 U2024 ( .A1(n1770), .A2(n1803), .B1(n1858), .B2(n1769), .ZN(n746)
         );
  AOI22_X1 U2025 ( .A1(n1770), .A2(n1804), .B1(n1859), .B2(n1769), .ZN(n745)
         );
  AOI22_X1 U2026 ( .A1(n1770), .A2(n1805), .B1(n1860), .B2(n1769), .ZN(n744)
         );
  AOI22_X1 U2027 ( .A1(n1770), .A2(n1806), .B1(n1861), .B2(n1769), .ZN(n743)
         );
  AOI22_X1 U2028 ( .A1(n1770), .A2(n1807), .B1(n1862), .B2(n1769), .ZN(n742)
         );
  AOI22_X1 U2029 ( .A1(n1770), .A2(n1809), .B1(n1863), .B2(n1769), .ZN(n741)
         );
  NOR2_X2 U2030 ( .A1(n1776), .A2(n1782), .ZN(n1772) );
  AOI22_X1 U2031 ( .A1(n1772), .A2(n1793), .B1(n1875), .B2(n1771), .ZN(n740)
         );
  AOI22_X1 U2032 ( .A1(n1772), .A2(n1794), .B1(n1876), .B2(n1771), .ZN(n739)
         );
  AOI22_X1 U2033 ( .A1(n1772), .A2(n1795), .B1(n1877), .B2(n1771), .ZN(n738)
         );
  AOI22_X1 U2034 ( .A1(n1772), .A2(n1796), .B1(n1878), .B2(n1771), .ZN(n737)
         );
  AOI22_X1 U2035 ( .A1(n1772), .A2(n1797), .B1(n1879), .B2(n1771), .ZN(n736)
         );
  AOI22_X1 U2036 ( .A1(n1772), .A2(n1798), .B1(n1880), .B2(n1771), .ZN(n735)
         );
  AOI22_X1 U2037 ( .A1(n1772), .A2(n1799), .B1(n1881), .B2(n1771), .ZN(n734)
         );
  AOI22_X1 U2038 ( .A1(n1772), .A2(n1800), .B1(n1882), .B2(n1771), .ZN(n733)
         );
  AOI22_X1 U2039 ( .A1(n1772), .A2(n1801), .B1(n1883), .B2(n1771), .ZN(n732)
         );
  AOI22_X1 U2040 ( .A1(n1772), .A2(n1802), .B1(n1884), .B2(n1771), .ZN(n731)
         );
  AOI22_X1 U2041 ( .A1(n1772), .A2(n1803), .B1(n1885), .B2(n1771), .ZN(n730)
         );
  AOI22_X1 U2042 ( .A1(n1772), .A2(n1804), .B1(n1886), .B2(n1771), .ZN(n729)
         );
  AOI22_X1 U2043 ( .A1(n1772), .A2(n1805), .B1(n1887), .B2(n1771), .ZN(n728)
         );
  AOI22_X1 U2044 ( .A1(n1772), .A2(n1806), .B1(n1888), .B2(n1771), .ZN(n727)
         );
  AOI22_X1 U2045 ( .A1(n1772), .A2(n1807), .B1(n1889), .B2(n1771), .ZN(n726)
         );
  AOI22_X1 U2046 ( .A1(n1772), .A2(n1809), .B1(n1890), .B2(n1771), .ZN(n725)
         );
  AOI22_X1 U2047 ( .A1(n1775), .A2(n1793), .B1(n1891), .B2(n1774), .ZN(n724)
         );
  AOI22_X1 U2048 ( .A1(n1775), .A2(n1794), .B1(n1892), .B2(n1774), .ZN(n723)
         );
  AOI22_X1 U2049 ( .A1(n1775), .A2(n1795), .B1(n1893), .B2(n1774), .ZN(n722)
         );
  AOI22_X1 U2050 ( .A1(n1775), .A2(n1796), .B1(n1894), .B2(n1774), .ZN(n721)
         );
  AOI22_X1 U2051 ( .A1(n1775), .A2(n1797), .B1(n1895), .B2(n1774), .ZN(n720)
         );
  AOI22_X1 U2052 ( .A1(n1775), .A2(n1798), .B1(n1896), .B2(n1774), .ZN(n719)
         );
  AOI22_X1 U2053 ( .A1(n1775), .A2(n1799), .B1(n1897), .B2(n1774), .ZN(n718)
         );
  AOI22_X1 U2054 ( .A1(n1775), .A2(n1800), .B1(n1898), .B2(n1774), .ZN(n717)
         );
  AOI22_X1 U2055 ( .A1(n1775), .A2(n1801), .B1(n1899), .B2(n1774), .ZN(n716)
         );
  AOI22_X1 U2056 ( .A1(n1775), .A2(n1802), .B1(n1900), .B2(n1774), .ZN(n715)
         );
  AOI22_X1 U2057 ( .A1(n1775), .A2(n1803), .B1(n1901), .B2(n1774), .ZN(n714)
         );
  AOI22_X1 U2058 ( .A1(n1775), .A2(n1804), .B1(n1902), .B2(n1774), .ZN(n713)
         );
  AOI22_X1 U2059 ( .A1(n1775), .A2(n1805), .B1(n1903), .B2(n1774), .ZN(n712)
         );
  AOI22_X1 U2060 ( .A1(n1775), .A2(n1806), .B1(n1904), .B2(n1774), .ZN(n711)
         );
  AOI22_X1 U2061 ( .A1(n1775), .A2(n1807), .B1(n1905), .B2(n1774), .ZN(n710)
         );
  AOI22_X1 U2062 ( .A1(n1775), .A2(n1809), .B1(n1906), .B2(n1774), .ZN(n709)
         );
  NOR2_X2 U2063 ( .A1(n1776), .A2(n1789), .ZN(n1778) );
  AOI22_X1 U2064 ( .A1(n1778), .A2(n1793), .B1(n1907), .B2(n1777), .ZN(n708)
         );
  AOI22_X1 U2065 ( .A1(n1778), .A2(n1794), .B1(n1908), .B2(n1777), .ZN(n707)
         );
  AOI22_X1 U2066 ( .A1(n1778), .A2(n1795), .B1(n1909), .B2(n1777), .ZN(n706)
         );
  AOI22_X1 U2067 ( .A1(n1778), .A2(n1796), .B1(n1910), .B2(n1777), .ZN(n705)
         );
  AOI22_X1 U2068 ( .A1(n1778), .A2(n1797), .B1(n1911), .B2(n1777), .ZN(n704)
         );
  AOI22_X1 U2069 ( .A1(n1778), .A2(n1798), .B1(n1912), .B2(n1777), .ZN(n703)
         );
  AOI22_X1 U2070 ( .A1(n1778), .A2(n1799), .B1(n1913), .B2(n1777), .ZN(n702)
         );
  AOI22_X1 U2071 ( .A1(n1778), .A2(n1800), .B1(n1914), .B2(n1777), .ZN(n701)
         );
  AOI22_X1 U2072 ( .A1(n1778), .A2(n1801), .B1(n1915), .B2(n1777), .ZN(n700)
         );
  AOI22_X1 U2073 ( .A1(n1778), .A2(n1802), .B1(n1916), .B2(n1777), .ZN(n699)
         );
  AOI22_X1 U2074 ( .A1(n1778), .A2(n1803), .B1(n1917), .B2(n1777), .ZN(n698)
         );
  AOI22_X1 U2075 ( .A1(n1778), .A2(n1804), .B1(n1918), .B2(n1777), .ZN(n697)
         );
  AOI22_X1 U2076 ( .A1(n1778), .A2(n1805), .B1(n1919), .B2(n1777), .ZN(n696)
         );
  AOI22_X1 U2077 ( .A1(n1778), .A2(n1806), .B1(n1920), .B2(n1777), .ZN(n695)
         );
  AOI22_X1 U2078 ( .A1(n1778), .A2(n1807), .B1(n1921), .B2(n1777), .ZN(n694)
         );
  AOI22_X1 U2079 ( .A1(n1778), .A2(n1809), .B1(n1922), .B2(n1777), .ZN(n693)
         );
  AOI22_X1 U2080 ( .A1(n1781), .A2(n1793), .B1(n1923), .B2(n1780), .ZN(n692)
         );
  AOI22_X1 U2081 ( .A1(n1781), .A2(n1794), .B1(n1924), .B2(n1780), .ZN(n691)
         );
  AOI22_X1 U2082 ( .A1(n1781), .A2(n1795), .B1(n1925), .B2(n1780), .ZN(n690)
         );
  AOI22_X1 U2083 ( .A1(n1781), .A2(n1796), .B1(n1926), .B2(n1780), .ZN(n689)
         );
  AOI22_X1 U2084 ( .A1(n1781), .A2(n1797), .B1(n1927), .B2(n1780), .ZN(n688)
         );
  AOI22_X1 U2085 ( .A1(n1781), .A2(n1798), .B1(n1928), .B2(n1780), .ZN(n687)
         );
  AOI22_X1 U2086 ( .A1(n1781), .A2(n1799), .B1(n1929), .B2(n1780), .ZN(n686)
         );
  AOI22_X1 U2087 ( .A1(n1781), .A2(n1800), .B1(n1930), .B2(n1780), .ZN(n685)
         );
  AOI22_X1 U2088 ( .A1(n1781), .A2(n1801), .B1(n1931), .B2(n1780), .ZN(n684)
         );
  AOI22_X1 U2089 ( .A1(n1781), .A2(n1802), .B1(n1932), .B2(n1780), .ZN(n683)
         );
  AOI22_X1 U2090 ( .A1(n1781), .A2(n1803), .B1(n1933), .B2(n1780), .ZN(n682)
         );
  AOI22_X1 U2091 ( .A1(n1781), .A2(n1804), .B1(n1934), .B2(n1780), .ZN(n681)
         );
  AOI22_X1 U2092 ( .A1(n1781), .A2(n1805), .B1(n1935), .B2(n1780), .ZN(n680)
         );
  AOI22_X1 U2093 ( .A1(n1781), .A2(n1806), .B1(n1936), .B2(n1780), .ZN(n679)
         );
  AOI22_X1 U2094 ( .A1(n1781), .A2(n1807), .B1(n1937), .B2(n1780), .ZN(n678)
         );
  AOI22_X1 U2095 ( .A1(n1781), .A2(n1809), .B1(n1938), .B2(n1780), .ZN(n677)
         );
  NOR2_X2 U2096 ( .A1(n1790), .A2(n1782), .ZN(n1784) );
  AOI22_X1 U2097 ( .A1(n1784), .A2(n1793), .B1(n2084), .B2(n1783), .ZN(n676)
         );
  AOI22_X1 U2098 ( .A1(n1784), .A2(n1794), .B1(n2085), .B2(n1783), .ZN(n675)
         );
  AOI22_X1 U2099 ( .A1(n1784), .A2(n1795), .B1(n2086), .B2(n1783), .ZN(n674)
         );
  AOI22_X1 U2100 ( .A1(n1784), .A2(n1796), .B1(n2087), .B2(n1783), .ZN(n673)
         );
  AOI22_X1 U2101 ( .A1(n1784), .A2(n1797), .B1(n2088), .B2(n1783), .ZN(n672)
         );
  AOI22_X1 U2102 ( .A1(n1784), .A2(n1798), .B1(n2089), .B2(n1783), .ZN(n671)
         );
  AOI22_X1 U2103 ( .A1(n1784), .A2(n1799), .B1(n2090), .B2(n1783), .ZN(n670)
         );
  AOI22_X1 U2104 ( .A1(n1784), .A2(n1800), .B1(n2091), .B2(n1783), .ZN(n669)
         );
  AOI22_X1 U2105 ( .A1(n1784), .A2(n1801), .B1(n2092), .B2(n1783), .ZN(n668)
         );
  AOI22_X1 U2106 ( .A1(n1784), .A2(n1802), .B1(n2093), .B2(n1783), .ZN(n667)
         );
  AOI22_X1 U2107 ( .A1(n1784), .A2(n1803), .B1(n2094), .B2(n1783), .ZN(n666)
         );
  AOI22_X1 U2108 ( .A1(n1784), .A2(n1804), .B1(n2095), .B2(n1783), .ZN(n665)
         );
  AOI22_X1 U2109 ( .A1(n1784), .A2(n1805), .B1(n2096), .B2(n1783), .ZN(n664)
         );
  AOI22_X1 U2110 ( .A1(n1784), .A2(n1806), .B1(n2097), .B2(n1783), .ZN(n663)
         );
  AOI22_X1 U2111 ( .A1(n1784), .A2(n1807), .B1(n2098), .B2(n1783), .ZN(n662)
         );
  AOI22_X1 U2112 ( .A1(n1784), .A2(n1809), .B1(n2099), .B2(n1783), .ZN(n661)
         );
  AOI22_X1 U2113 ( .A1(n1788), .A2(n1793), .B1(n2003), .B2(n1787), .ZN(n660)
         );
  AOI22_X1 U2114 ( .A1(n1788), .A2(n1794), .B1(n2004), .B2(n1787), .ZN(n659)
         );
  AOI22_X1 U2115 ( .A1(n1788), .A2(n1795), .B1(n2005), .B2(n1787), .ZN(n658)
         );
  AOI22_X1 U2116 ( .A1(n1788), .A2(n1796), .B1(n2006), .B2(n1787), .ZN(n657)
         );
  AOI22_X1 U2117 ( .A1(n1788), .A2(n1797), .B1(n2007), .B2(n1787), .ZN(n656)
         );
  AOI22_X1 U2118 ( .A1(n1788), .A2(n1798), .B1(n2008), .B2(n1787), .ZN(n655)
         );
  AOI22_X1 U2119 ( .A1(n1788), .A2(n1799), .B1(n2009), .B2(n1787), .ZN(n654)
         );
  AOI22_X1 U2120 ( .A1(n1788), .A2(n1800), .B1(n2010), .B2(n1787), .ZN(n653)
         );
  AOI22_X1 U2121 ( .A1(n1788), .A2(n1801), .B1(n2011), .B2(n1787), .ZN(n652)
         );
  AOI22_X1 U2122 ( .A1(n1788), .A2(n1802), .B1(n2012), .B2(n1787), .ZN(n651)
         );
  AOI22_X1 U2123 ( .A1(n1788), .A2(n1803), .B1(n2013), .B2(n1787), .ZN(n650)
         );
  AOI22_X1 U2124 ( .A1(n1788), .A2(n1804), .B1(n2014), .B2(n1787), .ZN(n649)
         );
  AOI22_X1 U2125 ( .A1(n1788), .A2(n1805), .B1(n2015), .B2(n1787), .ZN(n648)
         );
  AOI22_X1 U2126 ( .A1(n1788), .A2(n1806), .B1(n2016), .B2(n1787), .ZN(n647)
         );
  AOI22_X1 U2127 ( .A1(n1788), .A2(n1807), .B1(n2017), .B2(n1787), .ZN(n646)
         );
  AOI22_X1 U2128 ( .A1(n1788), .A2(n1809), .B1(n2018), .B2(n1787), .ZN(n645)
         );
  NOR2_X2 U2129 ( .A1(n1790), .A2(n1789), .ZN(n1792) );
  AOI22_X1 U2130 ( .A1(n1792), .A2(n1793), .B1(n2100), .B2(n1791), .ZN(n644)
         );
  AOI22_X1 U2131 ( .A1(n1792), .A2(n1794), .B1(n2101), .B2(n1791), .ZN(n643)
         );
  AOI22_X1 U2132 ( .A1(n1792), .A2(n1795), .B1(n2102), .B2(n1791), .ZN(n642)
         );
  AOI22_X1 U2133 ( .A1(n1792), .A2(n1796), .B1(n2103), .B2(n1791), .ZN(n641)
         );
  AOI22_X1 U2134 ( .A1(n1792), .A2(n1797), .B1(n2104), .B2(n1791), .ZN(n640)
         );
  AOI22_X1 U2135 ( .A1(n1792), .A2(n1798), .B1(n2105), .B2(n1791), .ZN(n639)
         );
  AOI22_X1 U2136 ( .A1(n1792), .A2(n1799), .B1(n2106), .B2(n1791), .ZN(n638)
         );
  AOI22_X1 U2137 ( .A1(n1792), .A2(n1800), .B1(n2107), .B2(n1791), .ZN(n637)
         );
  AOI22_X1 U2138 ( .A1(n1792), .A2(n1801), .B1(n2108), .B2(n1791), .ZN(n636)
         );
  AOI22_X1 U2139 ( .A1(n1792), .A2(n1802), .B1(n2109), .B2(n1791), .ZN(n635)
         );
  AOI22_X1 U2140 ( .A1(n1792), .A2(n1803), .B1(n2110), .B2(n1791), .ZN(n634)
         );
  AOI22_X1 U2141 ( .A1(n1792), .A2(n1804), .B1(n2111), .B2(n1791), .ZN(n633)
         );
  AOI22_X1 U2142 ( .A1(n1792), .A2(n1805), .B1(n2112), .B2(n1791), .ZN(n632)
         );
  AOI22_X1 U2143 ( .A1(n1792), .A2(n1806), .B1(n2113), .B2(n1791), .ZN(n631)
         );
  AOI22_X1 U2144 ( .A1(n1792), .A2(n1807), .B1(n2114), .B2(n1791), .ZN(n630)
         );
  AOI22_X1 U2145 ( .A1(n1792), .A2(n1809), .B1(n2115), .B2(n1791), .ZN(n629)
         );
  AOI22_X1 U2146 ( .A1(n1810), .A2(n1793), .B1(n2019), .B2(n1808), .ZN(n628)
         );
  AOI22_X1 U2147 ( .A1(n1810), .A2(n1794), .B1(n2020), .B2(n1808), .ZN(n627)
         );
  AOI22_X1 U2148 ( .A1(n1810), .A2(n1795), .B1(n2021), .B2(n1808), .ZN(n626)
         );
  AOI22_X1 U2149 ( .A1(n1810), .A2(n1796), .B1(n2022), .B2(n1808), .ZN(n625)
         );
  AOI22_X1 U2150 ( .A1(n1810), .A2(n1797), .B1(n2023), .B2(n1808), .ZN(n624)
         );
  AOI22_X1 U2151 ( .A1(n1810), .A2(n1798), .B1(n2024), .B2(n1808), .ZN(n623)
         );
  AOI22_X1 U2152 ( .A1(n1810), .A2(n1799), .B1(n2025), .B2(n1808), .ZN(n622)
         );
  AOI22_X1 U2153 ( .A1(n1810), .A2(n1800), .B1(n2026), .B2(n1808), .ZN(n621)
         );
  AOI22_X1 U2154 ( .A1(n1810), .A2(n1801), .B1(n2027), .B2(n1808), .ZN(n620)
         );
  AOI22_X1 U2155 ( .A1(n1810), .A2(n1802), .B1(n2028), .B2(n1808), .ZN(n619)
         );
  AOI22_X1 U2156 ( .A1(n1810), .A2(n1803), .B1(n2029), .B2(n1808), .ZN(n618)
         );
  AOI22_X1 U2157 ( .A1(n1810), .A2(n1804), .B1(n2030), .B2(n1808), .ZN(n617)
         );
  AOI22_X1 U2158 ( .A1(n1810), .A2(n1805), .B1(n2031), .B2(n1808), .ZN(n616)
         );
  AOI22_X1 U2159 ( .A1(n1810), .A2(n1806), .B1(n2032), .B2(n1808), .ZN(n615)
         );
  AOI22_X1 U2160 ( .A1(n1810), .A2(n1807), .B1(n2033), .B2(n1808), .ZN(n614)
         );
  AOI22_X1 U2161 ( .A1(n1810), .A2(n1809), .B1(n2034), .B2(n1808), .ZN(n613)
         );
  NAND3_X1 U2162 ( .A1(\ctrl_conv_output_inst/m_pre_valid_y ), .A2(n1812), 
        .A3(n1811), .ZN(n1813) );
  OAI21_X1 U2163 ( .B1(n1814), .B2(n1836), .A(n1813), .ZN(n612) );
endmodule

