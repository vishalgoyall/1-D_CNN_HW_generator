
module conv_30_9_11_1 ( clk, reset, s_data_in_x, s_valid_x, s_ready_x, 
        m_data_out_y, m_valid_y, m_ready_y );
  input [10:0] s_data_in_x;
  output [10:0] m_data_out_y;
  input clk, reset, s_valid_x, m_ready_y;
  output s_ready_x, m_valid_y;
  wire   conv_done, N29, \xmem_inst/N24 , \xmem_inst/N22 , \xmem_inst/N19 ,
         \xmem_inst/N18 , \xmem_inst/N16 , \xmem_inst/mem[29][10] ,
         \xmem_inst/mem[29][9] , \xmem_inst/mem[29][8] ,
         \xmem_inst/mem[29][7] , \xmem_inst/mem[29][6] ,
         \xmem_inst/mem[29][5] , \xmem_inst/mem[29][4] ,
         \xmem_inst/mem[29][3] , \xmem_inst/mem[29][2] ,
         \xmem_inst/mem[29][1] , \xmem_inst/mem[29][0] ,
         \xmem_inst/mem[28][10] , \xmem_inst/mem[28][9] ,
         \xmem_inst/mem[28][8] , \xmem_inst/mem[28][7] ,
         \xmem_inst/mem[28][6] , \xmem_inst/mem[28][5] ,
         \xmem_inst/mem[28][4] , \xmem_inst/mem[28][3] ,
         \xmem_inst/mem[28][2] , \xmem_inst/mem[28][1] ,
         \xmem_inst/mem[28][0] , \xmem_inst/mem[27][10] ,
         \xmem_inst/mem[27][9] , \xmem_inst/mem[27][8] ,
         \xmem_inst/mem[27][7] , \xmem_inst/mem[27][6] ,
         \xmem_inst/mem[27][5] , \xmem_inst/mem[27][4] ,
         \xmem_inst/mem[27][3] , \xmem_inst/mem[27][2] ,
         \xmem_inst/mem[27][1] , \xmem_inst/mem[27][0] ,
         \xmem_inst/mem[26][10] , \xmem_inst/mem[26][9] ,
         \xmem_inst/mem[26][8] , \xmem_inst/mem[26][7] ,
         \xmem_inst/mem[26][6] , \xmem_inst/mem[26][5] ,
         \xmem_inst/mem[26][4] , \xmem_inst/mem[26][3] ,
         \xmem_inst/mem[26][2] , \xmem_inst/mem[26][1] ,
         \xmem_inst/mem[26][0] , \xmem_inst/mem[25][10] ,
         \xmem_inst/mem[25][9] , \xmem_inst/mem[25][8] ,
         \xmem_inst/mem[25][7] , \xmem_inst/mem[25][6] ,
         \xmem_inst/mem[25][5] , \xmem_inst/mem[25][4] ,
         \xmem_inst/mem[25][3] , \xmem_inst/mem[25][2] ,
         \xmem_inst/mem[25][1] , \xmem_inst/mem[25][0] ,
         \xmem_inst/mem[24][10] , \xmem_inst/mem[24][9] ,
         \xmem_inst/mem[24][8] , \xmem_inst/mem[24][7] ,
         \xmem_inst/mem[24][6] , \xmem_inst/mem[24][5] ,
         \xmem_inst/mem[24][4] , \xmem_inst/mem[24][3] ,
         \xmem_inst/mem[24][2] , \xmem_inst/mem[24][1] ,
         \xmem_inst/mem[24][0] , \xmem_inst/mem[23][10] ,
         \xmem_inst/mem[23][9] , \xmem_inst/mem[23][8] ,
         \xmem_inst/mem[23][7] , \xmem_inst/mem[23][6] ,
         \xmem_inst/mem[23][5] , \xmem_inst/mem[23][4] ,
         \xmem_inst/mem[23][3] , \xmem_inst/mem[23][2] ,
         \xmem_inst/mem[23][1] , \xmem_inst/mem[23][0] ,
         \xmem_inst/mem[22][10] , \xmem_inst/mem[22][9] ,
         \xmem_inst/mem[22][8] , \xmem_inst/mem[22][7] ,
         \xmem_inst/mem[22][6] , \xmem_inst/mem[22][5] ,
         \xmem_inst/mem[22][4] , \xmem_inst/mem[22][3] ,
         \xmem_inst/mem[22][2] , \xmem_inst/mem[22][1] ,
         \xmem_inst/mem[22][0] , \xmem_inst/mem[21][10] ,
         \xmem_inst/mem[21][9] , \xmem_inst/mem[21][8] ,
         \xmem_inst/mem[21][7] , \xmem_inst/mem[21][6] ,
         \xmem_inst/mem[21][5] , \xmem_inst/mem[21][4] ,
         \xmem_inst/mem[21][3] , \xmem_inst/mem[21][2] ,
         \xmem_inst/mem[21][1] , \xmem_inst/mem[21][0] ,
         \xmem_inst/mem[20][10] , \xmem_inst/mem[20][9] ,
         \xmem_inst/mem[20][8] , \xmem_inst/mem[20][7] ,
         \xmem_inst/mem[20][6] , \xmem_inst/mem[20][5] ,
         \xmem_inst/mem[20][4] , \xmem_inst/mem[20][3] ,
         \xmem_inst/mem[20][2] , \xmem_inst/mem[20][1] ,
         \xmem_inst/mem[20][0] , \xmem_inst/mem[19][10] ,
         \xmem_inst/mem[19][9] , \xmem_inst/mem[19][8] ,
         \xmem_inst/mem[19][7] , \xmem_inst/mem[19][6] ,
         \xmem_inst/mem[19][5] , \xmem_inst/mem[19][4] ,
         \xmem_inst/mem[19][3] , \xmem_inst/mem[19][2] ,
         \xmem_inst/mem[19][1] , \xmem_inst/mem[19][0] ,
         \xmem_inst/mem[18][10] , \xmem_inst/mem[18][9] ,
         \xmem_inst/mem[18][8] , \xmem_inst/mem[18][7] ,
         \xmem_inst/mem[18][6] , \xmem_inst/mem[18][5] ,
         \xmem_inst/mem[18][4] , \xmem_inst/mem[18][3] ,
         \xmem_inst/mem[18][2] , \xmem_inst/mem[18][1] ,
         \xmem_inst/mem[18][0] , \xmem_inst/mem[17][10] ,
         \xmem_inst/mem[17][9] , \xmem_inst/mem[17][8] ,
         \xmem_inst/mem[17][7] , \xmem_inst/mem[17][6] ,
         \xmem_inst/mem[17][5] , \xmem_inst/mem[17][4] ,
         \xmem_inst/mem[17][3] , \xmem_inst/mem[17][2] ,
         \xmem_inst/mem[17][1] , \xmem_inst/mem[17][0] ,
         \xmem_inst/mem[16][10] , \xmem_inst/mem[16][9] ,
         \xmem_inst/mem[16][8] , \xmem_inst/mem[16][7] ,
         \xmem_inst/mem[16][6] , \xmem_inst/mem[16][5] ,
         \xmem_inst/mem[16][4] , \xmem_inst/mem[16][3] ,
         \xmem_inst/mem[16][2] , \xmem_inst/mem[16][1] ,
         \xmem_inst/mem[16][0] , \xmem_inst/mem[15][10] ,
         \xmem_inst/mem[15][9] , \xmem_inst/mem[15][8] ,
         \xmem_inst/mem[15][7] , \xmem_inst/mem[15][6] ,
         \xmem_inst/mem[15][5] , \xmem_inst/mem[15][4] ,
         \xmem_inst/mem[15][3] , \xmem_inst/mem[15][2] ,
         \xmem_inst/mem[15][1] , \xmem_inst/mem[15][0] ,
         \xmem_inst/mem[14][10] , \xmem_inst/mem[14][9] ,
         \xmem_inst/mem[14][8] , \xmem_inst/mem[14][7] ,
         \xmem_inst/mem[14][6] , \xmem_inst/mem[14][5] ,
         \xmem_inst/mem[14][4] , \xmem_inst/mem[14][3] ,
         \xmem_inst/mem[14][2] , \xmem_inst/mem[14][1] ,
         \xmem_inst/mem[14][0] , \xmem_inst/mem[13][10] ,
         \xmem_inst/mem[13][9] , \xmem_inst/mem[13][8] ,
         \xmem_inst/mem[13][7] , \xmem_inst/mem[13][6] ,
         \xmem_inst/mem[13][5] , \xmem_inst/mem[13][4] ,
         \xmem_inst/mem[13][3] , \xmem_inst/mem[13][2] ,
         \xmem_inst/mem[13][1] , \xmem_inst/mem[13][0] ,
         \xmem_inst/mem[12][10] , \xmem_inst/mem[12][9] ,
         \xmem_inst/mem[12][8] , \xmem_inst/mem[12][7] ,
         \xmem_inst/mem[12][6] , \xmem_inst/mem[12][5] ,
         \xmem_inst/mem[12][4] , \xmem_inst/mem[12][3] ,
         \xmem_inst/mem[12][2] , \xmem_inst/mem[12][1] ,
         \xmem_inst/mem[12][0] , \xmem_inst/mem[11][10] ,
         \xmem_inst/mem[11][9] , \xmem_inst/mem[11][8] ,
         \xmem_inst/mem[11][7] , \xmem_inst/mem[11][6] ,
         \xmem_inst/mem[11][5] , \xmem_inst/mem[11][4] ,
         \xmem_inst/mem[11][3] , \xmem_inst/mem[11][2] ,
         \xmem_inst/mem[11][1] , \xmem_inst/mem[11][0] ,
         \xmem_inst/mem[10][10] , \xmem_inst/mem[10][9] ,
         \xmem_inst/mem[10][8] , \xmem_inst/mem[10][7] ,
         \xmem_inst/mem[10][6] , \xmem_inst/mem[10][5] ,
         \xmem_inst/mem[10][4] , \xmem_inst/mem[10][3] ,
         \xmem_inst/mem[10][2] , \xmem_inst/mem[10][1] ,
         \xmem_inst/mem[10][0] , \xmem_inst/mem[9][10] , \xmem_inst/mem[9][9] ,
         \xmem_inst/mem[9][8] , \xmem_inst/mem[9][7] , \xmem_inst/mem[9][6] ,
         \xmem_inst/mem[9][5] , \xmem_inst/mem[9][4] , \xmem_inst/mem[9][3] ,
         \xmem_inst/mem[9][2] , \xmem_inst/mem[9][1] , \xmem_inst/mem[9][0] ,
         \xmem_inst/mem[8][10] , \xmem_inst/mem[8][9] , \xmem_inst/mem[8][8] ,
         \xmem_inst/mem[8][7] , \xmem_inst/mem[8][6] , \xmem_inst/mem[8][5] ,
         \xmem_inst/mem[8][4] , \xmem_inst/mem[8][3] , \xmem_inst/mem[8][2] ,
         \xmem_inst/mem[8][1] , \xmem_inst/mem[8][0] , \xmem_inst/mem[7][10] ,
         \xmem_inst/mem[7][9] , \xmem_inst/mem[7][8] , \xmem_inst/mem[7][7] ,
         \xmem_inst/mem[7][6] , \xmem_inst/mem[7][5] , \xmem_inst/mem[7][4] ,
         \xmem_inst/mem[7][3] , \xmem_inst/mem[7][2] , \xmem_inst/mem[7][1] ,
         \xmem_inst/mem[7][0] , \xmem_inst/mem[6][10] , \xmem_inst/mem[6][9] ,
         \xmem_inst/mem[6][8] , \xmem_inst/mem[6][7] , \xmem_inst/mem[6][6] ,
         \xmem_inst/mem[6][5] , \xmem_inst/mem[6][4] , \xmem_inst/mem[6][3] ,
         \xmem_inst/mem[6][2] , \xmem_inst/mem[6][1] , \xmem_inst/mem[6][0] ,
         \xmem_inst/mem[5][10] , \xmem_inst/mem[5][9] , \xmem_inst/mem[5][8] ,
         \xmem_inst/mem[5][7] , \xmem_inst/mem[5][6] , \xmem_inst/mem[5][5] ,
         \xmem_inst/mem[5][4] , \xmem_inst/mem[5][3] , \xmem_inst/mem[5][2] ,
         \xmem_inst/mem[5][1] , \xmem_inst/mem[5][0] , \xmem_inst/mem[4][10] ,
         \xmem_inst/mem[4][9] , \xmem_inst/mem[4][8] , \xmem_inst/mem[4][7] ,
         \xmem_inst/mem[4][6] , \xmem_inst/mem[4][5] , \xmem_inst/mem[4][4] ,
         \xmem_inst/mem[4][3] , \xmem_inst/mem[4][2] , \xmem_inst/mem[4][1] ,
         \xmem_inst/mem[4][0] , \xmem_inst/mem[3][10] , \xmem_inst/mem[3][9] ,
         \xmem_inst/mem[3][8] , \xmem_inst/mem[3][7] , \xmem_inst/mem[3][6] ,
         \xmem_inst/mem[3][5] , \xmem_inst/mem[3][4] , \xmem_inst/mem[3][3] ,
         \xmem_inst/mem[3][2] , \xmem_inst/mem[3][1] , \xmem_inst/mem[3][0] ,
         \xmem_inst/mem[2][10] , \xmem_inst/mem[2][9] , \xmem_inst/mem[2][8] ,
         \xmem_inst/mem[2][7] , \xmem_inst/mem[2][6] , \xmem_inst/mem[2][5] ,
         \xmem_inst/mem[2][4] , \xmem_inst/mem[2][3] , \xmem_inst/mem[2][2] ,
         \xmem_inst/mem[2][1] , \xmem_inst/mem[2][0] , \xmem_inst/mem[1][10] ,
         \xmem_inst/mem[1][9] , \xmem_inst/mem[1][8] , \xmem_inst/mem[1][7] ,
         \xmem_inst/mem[1][6] , \xmem_inst/mem[1][5] , \xmem_inst/mem[1][4] ,
         \xmem_inst/mem[1][3] , \xmem_inst/mem[1][2] , \xmem_inst/mem[1][1] ,
         \xmem_inst/mem[1][0] , \xmem_inst/mem[0][10] , \xmem_inst/mem[0][9] ,
         \xmem_inst/mem[0][8] , \xmem_inst/mem[0][7] , \xmem_inst/mem[0][6] ,
         \xmem_inst/mem[0][5] , \xmem_inst/mem[0][4] , \xmem_inst/mem[0][3] ,
         \xmem_inst/mem[0][2] , \xmem_inst/mem[0][1] , \xmem_inst/mem[0][0] ,
         \ctrl_conv_output_inst/N77 , \ctrl_conv_output_inst/N74 ,
         \ctrl_conv_output_inst/m_pre_valid_y ,
         \ctrl_conv_output_inst/m_pre_pre_valid_y , n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1155, n1156, n1157, n1158,
         n1159, \DP_OP_65J1_122_2282/n664 , \DP_OP_65J1_122_2282/n663 , n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520;
  wire   [4:0] xmem_addr;
  wire   [10:0] xmem_data;
  wire   [3:0] fmem_addr;
  wire   [10:0] fmem_data;
  wire   [4:0] \ctrl_conv_output_inst/cnt_conv ;
  wire   [10:0] \mac_unit_inst/adder_reg ;
  wire   [10:0] \mac_unit_inst/x_mult_f_reg ;
  assign m_data_out_y[10] = 1'b0;

  DFF_X1 \xmem_inst/data_out_reg[2]  ( .D(\xmem_inst/N24 ), .CK(clk), .Q(
        xmem_data[2]), .QN(n2474) );
  DFF_X1 \xmem_inst/data_out_reg[4]  ( .D(\xmem_inst/N22 ), .CK(clk), .Q(n1218), .QN(n2482) );
  DFF_X1 \xmem_inst/data_out_reg[8]  ( .D(\xmem_inst/N18 ), .CK(clk), .QN(
        n2477) );
  DFF_X1 \ctrl_conv_output_inst/conv_done_reg  ( .D(
        \ctrl_conv_output_inst/N77 ), .CK(clk), .Q(conv_done) );
  DFF_X1 \ctrl_conv_output_inst/m_pre_pre_valid_y_reg  ( .D(n1159), .CK(clk), 
        .Q(\ctrl_conv_output_inst/m_pre_pre_valid_y ), .QN(n2490) );
  DFF_X1 \ctrl_conv_output_inst/m_pre_valid_y_reg  ( .D(n806), .CK(clk), .Q(
        \ctrl_conv_output_inst/m_pre_valid_y ), .QN(n2503) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[4]  ( .D(n1158), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [4]) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[0]  ( .D(n1157), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [0]), .QN(n2492) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[1]  ( .D(n1156), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [1]), .QN(n2497) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[2]  ( .D(n1155), .CK(clk), .Q(
        \ctrl_conv_output_inst/cnt_conv [2]), .QN(n2501) );
  DFF_X1 \ctrl_conv_output_inst/m_valid_y_reg  ( .D(n1153), .CK(clk), .Q(
        m_valid_y) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[4]  ( .D(n1147), .CK(clk), .Q(
        xmem_addr[4]) );
  DFF_X1 \ctrl_xmem_write_inst/s_ready_reg  ( .D(n1152), .CK(clk), .Q(
        s_ready_x), .QN(n2511) );
  DFF_X1 conv_pre_start_reg ( .D(N29), .CK(clk), .QN(n2512) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[0]  ( .D(n1151), .CK(clk), .Q(
        xmem_addr[0]), .QN(n2493) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[1]  ( .D(n1150), .CK(clk), .Q(
        xmem_addr[1]), .QN(n2502) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[2]  ( .D(n1149), .CK(clk), .Q(
        xmem_addr[2]) );
  DFF_X1 \xmem_inst/mem_reg[24][0]  ( .D(n882), .CK(clk), .Q(
        \xmem_inst/mem[24][0] ) );
  DFF_X1 \xmem_inst/mem_reg[24][1]  ( .D(n881), .CK(clk), .Q(
        \xmem_inst/mem[24][1] ) );
  DFF_X1 \xmem_inst/mem_reg[24][2]  ( .D(n880), .CK(clk), .Q(
        \xmem_inst/mem[24][2] ) );
  DFF_X1 \xmem_inst/mem_reg[24][3]  ( .D(n879), .CK(clk), .Q(
        \xmem_inst/mem[24][3] ) );
  DFF_X1 \xmem_inst/mem_reg[24][4]  ( .D(n878), .CK(clk), .Q(
        \xmem_inst/mem[24][4] ) );
  DFF_X1 \xmem_inst/mem_reg[24][5]  ( .D(n877), .CK(clk), .Q(
        \xmem_inst/mem[24][5] ) );
  DFF_X1 \xmem_inst/mem_reg[24][6]  ( .D(n876), .CK(clk), .Q(
        \xmem_inst/mem[24][6] ) );
  DFF_X1 \xmem_inst/mem_reg[24][7]  ( .D(n875), .CK(clk), .Q(
        \xmem_inst/mem[24][7] ) );
  DFF_X1 \xmem_inst/mem_reg[24][8]  ( .D(n874), .CK(clk), .Q(
        \xmem_inst/mem[24][8] ) );
  DFF_X1 \xmem_inst/mem_reg[24][9]  ( .D(n873), .CK(clk), .Q(
        \xmem_inst/mem[24][9] ) );
  DFF_X1 \xmem_inst/mem_reg[24][10]  ( .D(n872), .CK(clk), .Q(
        \xmem_inst/mem[24][10] ) );
  DFF_X1 \xmem_inst/mem_reg[25][0]  ( .D(n871), .CK(clk), .Q(
        \xmem_inst/mem[25][0] ) );
  DFF_X1 \xmem_inst/mem_reg[25][1]  ( .D(n870), .CK(clk), .Q(
        \xmem_inst/mem[25][1] ) );
  DFF_X1 \xmem_inst/mem_reg[25][2]  ( .D(n869), .CK(clk), .Q(
        \xmem_inst/mem[25][2] ) );
  DFF_X1 \xmem_inst/mem_reg[25][3]  ( .D(n868), .CK(clk), .Q(
        \xmem_inst/mem[25][3] ) );
  DFF_X1 \xmem_inst/mem_reg[25][4]  ( .D(n867), .CK(clk), .Q(
        \xmem_inst/mem[25][4] ) );
  DFF_X1 \xmem_inst/mem_reg[25][5]  ( .D(n866), .CK(clk), .Q(
        \xmem_inst/mem[25][5] ) );
  DFF_X1 \xmem_inst/mem_reg[25][6]  ( .D(n865), .CK(clk), .Q(
        \xmem_inst/mem[25][6] ) );
  DFF_X1 \xmem_inst/mem_reg[25][7]  ( .D(n864), .CK(clk), .Q(
        \xmem_inst/mem[25][7] ) );
  DFF_X1 \xmem_inst/mem_reg[25][8]  ( .D(n863), .CK(clk), .Q(
        \xmem_inst/mem[25][8] ) );
  DFF_X1 \xmem_inst/mem_reg[25][9]  ( .D(n862), .CK(clk), .Q(
        \xmem_inst/mem[25][9] ) );
  DFF_X1 \xmem_inst/mem_reg[25][10]  ( .D(n861), .CK(clk), .Q(
        \xmem_inst/mem[25][10] ) );
  DFF_X1 \xmem_inst/mem_reg[26][0]  ( .D(n860), .CK(clk), .Q(
        \xmem_inst/mem[26][0] ) );
  DFF_X1 \xmem_inst/mem_reg[26][1]  ( .D(n859), .CK(clk), .Q(
        \xmem_inst/mem[26][1] ) );
  DFF_X1 \xmem_inst/mem_reg[26][2]  ( .D(n858), .CK(clk), .Q(
        \xmem_inst/mem[26][2] ) );
  DFF_X1 \xmem_inst/mem_reg[26][3]  ( .D(n857), .CK(clk), .Q(
        \xmem_inst/mem[26][3] ) );
  DFF_X1 \xmem_inst/mem_reg[26][4]  ( .D(n856), .CK(clk), .Q(
        \xmem_inst/mem[26][4] ) );
  DFF_X1 \xmem_inst/mem_reg[26][5]  ( .D(n855), .CK(clk), .Q(
        \xmem_inst/mem[26][5] ) );
  DFF_X1 \xmem_inst/mem_reg[26][6]  ( .D(n854), .CK(clk), .Q(
        \xmem_inst/mem[26][6] ) );
  DFF_X1 \xmem_inst/mem_reg[26][7]  ( .D(n853), .CK(clk), .Q(
        \xmem_inst/mem[26][7] ) );
  DFF_X1 \xmem_inst/mem_reg[26][8]  ( .D(n852), .CK(clk), .Q(
        \xmem_inst/mem[26][8] ) );
  DFF_X1 \xmem_inst/mem_reg[26][9]  ( .D(n851), .CK(clk), .Q(
        \xmem_inst/mem[26][9] ) );
  DFF_X1 \xmem_inst/mem_reg[26][10]  ( .D(n850), .CK(clk), .Q(
        \xmem_inst/mem[26][10] ) );
  DFF_X1 \xmem_inst/mem_reg[27][0]  ( .D(n849), .CK(clk), .Q(
        \xmem_inst/mem[27][0] ) );
  DFF_X1 \xmem_inst/mem_reg[27][1]  ( .D(n848), .CK(clk), .Q(
        \xmem_inst/mem[27][1] ) );
  DFF_X1 \xmem_inst/mem_reg[27][2]  ( .D(n847), .CK(clk), .Q(
        \xmem_inst/mem[27][2] ) );
  DFF_X1 \xmem_inst/mem_reg[27][3]  ( .D(n846), .CK(clk), .Q(
        \xmem_inst/mem[27][3] ) );
  DFF_X1 \xmem_inst/mem_reg[27][4]  ( .D(n845), .CK(clk), .Q(
        \xmem_inst/mem[27][4] ) );
  DFF_X1 \xmem_inst/mem_reg[27][5]  ( .D(n844), .CK(clk), .Q(
        \xmem_inst/mem[27][5] ) );
  DFF_X1 \xmem_inst/mem_reg[27][6]  ( .D(n843), .CK(clk), .Q(
        \xmem_inst/mem[27][6] ) );
  DFF_X1 \xmem_inst/mem_reg[27][7]  ( .D(n842), .CK(clk), .Q(
        \xmem_inst/mem[27][7] ) );
  DFF_X1 \xmem_inst/mem_reg[27][8]  ( .D(n841), .CK(clk), .Q(
        \xmem_inst/mem[27][8] ) );
  DFF_X1 \xmem_inst/mem_reg[27][9]  ( .D(n840), .CK(clk), .Q(
        \xmem_inst/mem[27][9] ) );
  DFF_X1 \xmem_inst/mem_reg[27][10]  ( .D(n839), .CK(clk), .Q(
        \xmem_inst/mem[27][10] ) );
  DFF_X1 \xmem_inst/mem_reg[28][0]  ( .D(n838), .CK(clk), .Q(
        \xmem_inst/mem[28][0] ) );
  DFF_X1 \xmem_inst/mem_reg[28][1]  ( .D(n837), .CK(clk), .Q(
        \xmem_inst/mem[28][1] ) );
  DFF_X1 \xmem_inst/mem_reg[28][2]  ( .D(n836), .CK(clk), .Q(
        \xmem_inst/mem[28][2] ) );
  DFF_X1 \xmem_inst/mem_reg[28][3]  ( .D(n835), .CK(clk), .Q(
        \xmem_inst/mem[28][3] ) );
  DFF_X1 \xmem_inst/mem_reg[28][4]  ( .D(n834), .CK(clk), .Q(
        \xmem_inst/mem[28][4] ) );
  DFF_X1 \xmem_inst/mem_reg[28][5]  ( .D(n833), .CK(clk), .Q(
        \xmem_inst/mem[28][5] ) );
  DFF_X1 \xmem_inst/mem_reg[28][6]  ( .D(n832), .CK(clk), .Q(
        \xmem_inst/mem[28][6] ) );
  DFF_X1 \xmem_inst/mem_reg[28][7]  ( .D(n831), .CK(clk), .Q(
        \xmem_inst/mem[28][7] ) );
  DFF_X1 \xmem_inst/mem_reg[28][8]  ( .D(n830), .CK(clk), .Q(
        \xmem_inst/mem[28][8] ) );
  DFF_X1 \xmem_inst/mem_reg[28][9]  ( .D(n829), .CK(clk), .Q(
        \xmem_inst/mem[28][9] ) );
  DFF_X1 \xmem_inst/mem_reg[28][10]  ( .D(n828), .CK(clk), .Q(
        \xmem_inst/mem[28][10] ) );
  DFF_X1 \ctrl_xmem_write_inst/mem_addr_reg[3]  ( .D(n1148), .CK(clk), .Q(
        xmem_addr[3]), .QN(n2495) );
  DFF_X1 \xmem_inst/mem_reg[8][0]  ( .D(n1058), .CK(clk), .Q(
        \xmem_inst/mem[8][0] ) );
  DFF_X1 \xmem_inst/mem_reg[8][1]  ( .D(n1057), .CK(clk), .Q(
        \xmem_inst/mem[8][1] ) );
  DFF_X1 \xmem_inst/mem_reg[8][2]  ( .D(n1056), .CK(clk), .Q(
        \xmem_inst/mem[8][2] ) );
  DFF_X1 \xmem_inst/mem_reg[8][3]  ( .D(n1055), .CK(clk), .Q(
        \xmem_inst/mem[8][3] ) );
  DFF_X1 \xmem_inst/mem_reg[8][4]  ( .D(n1054), .CK(clk), .Q(
        \xmem_inst/mem[8][4] ) );
  DFF_X1 \xmem_inst/mem_reg[8][5]  ( .D(n1053), .CK(clk), .Q(
        \xmem_inst/mem[8][5] ) );
  DFF_X1 \xmem_inst/mem_reg[8][6]  ( .D(n1052), .CK(clk), .Q(
        \xmem_inst/mem[8][6] ) );
  DFF_X1 \xmem_inst/mem_reg[8][7]  ( .D(n1051), .CK(clk), .Q(
        \xmem_inst/mem[8][7] ) );
  DFF_X1 \xmem_inst/mem_reg[8][8]  ( .D(n1050), .CK(clk), .Q(
        \xmem_inst/mem[8][8] ) );
  DFF_X1 \xmem_inst/mem_reg[8][9]  ( .D(n1049), .CK(clk), .Q(
        \xmem_inst/mem[8][9] ) );
  DFF_X1 \xmem_inst/mem_reg[8][10]  ( .D(n1048), .CK(clk), .Q(
        \xmem_inst/mem[8][10] ) );
  DFF_X1 \xmem_inst/mem_reg[9][0]  ( .D(n1047), .CK(clk), .Q(
        \xmem_inst/mem[9][0] ) );
  DFF_X1 \xmem_inst/mem_reg[9][1]  ( .D(n1046), .CK(clk), .Q(
        \xmem_inst/mem[9][1] ) );
  DFF_X1 \xmem_inst/mem_reg[9][2]  ( .D(n1045), .CK(clk), .Q(
        \xmem_inst/mem[9][2] ) );
  DFF_X1 \xmem_inst/mem_reg[9][3]  ( .D(n1044), .CK(clk), .Q(
        \xmem_inst/mem[9][3] ) );
  DFF_X1 \xmem_inst/mem_reg[9][4]  ( .D(n1043), .CK(clk), .Q(
        \xmem_inst/mem[9][4] ) );
  DFF_X1 \xmem_inst/mem_reg[9][5]  ( .D(n1042), .CK(clk), .Q(
        \xmem_inst/mem[9][5] ) );
  DFF_X1 \xmem_inst/mem_reg[9][6]  ( .D(n1041), .CK(clk), .Q(
        \xmem_inst/mem[9][6] ) );
  DFF_X1 \xmem_inst/mem_reg[9][7]  ( .D(n1040), .CK(clk), .Q(
        \xmem_inst/mem[9][7] ) );
  DFF_X1 \xmem_inst/mem_reg[9][8]  ( .D(n1039), .CK(clk), .Q(
        \xmem_inst/mem[9][8] ) );
  DFF_X1 \xmem_inst/mem_reg[9][9]  ( .D(n1038), .CK(clk), .Q(
        \xmem_inst/mem[9][9] ) );
  DFF_X1 \xmem_inst/mem_reg[9][10]  ( .D(n1037), .CK(clk), .Q(
        \xmem_inst/mem[9][10] ) );
  DFF_X1 \xmem_inst/mem_reg[10][0]  ( .D(n1036), .CK(clk), .Q(
        \xmem_inst/mem[10][0] ) );
  DFF_X1 \xmem_inst/mem_reg[10][1]  ( .D(n1035), .CK(clk), .Q(
        \xmem_inst/mem[10][1] ) );
  DFF_X1 \xmem_inst/mem_reg[10][2]  ( .D(n1034), .CK(clk), .Q(
        \xmem_inst/mem[10][2] ) );
  DFF_X1 \xmem_inst/mem_reg[10][3]  ( .D(n1033), .CK(clk), .Q(
        \xmem_inst/mem[10][3] ) );
  DFF_X1 \xmem_inst/mem_reg[10][4]  ( .D(n1032), .CK(clk), .Q(
        \xmem_inst/mem[10][4] ) );
  DFF_X1 \xmem_inst/mem_reg[10][5]  ( .D(n1031), .CK(clk), .Q(
        \xmem_inst/mem[10][5] ) );
  DFF_X1 \xmem_inst/mem_reg[10][6]  ( .D(n1030), .CK(clk), .Q(
        \xmem_inst/mem[10][6] ) );
  DFF_X1 \xmem_inst/mem_reg[10][7]  ( .D(n1029), .CK(clk), .Q(
        \xmem_inst/mem[10][7] ) );
  DFF_X1 \xmem_inst/mem_reg[10][8]  ( .D(n1028), .CK(clk), .Q(
        \xmem_inst/mem[10][8] ) );
  DFF_X1 \xmem_inst/mem_reg[10][9]  ( .D(n1027), .CK(clk), .Q(
        \xmem_inst/mem[10][9] ) );
  DFF_X1 \xmem_inst/mem_reg[10][10]  ( .D(n1026), .CK(clk), .Q(
        \xmem_inst/mem[10][10] ) );
  DFF_X1 \xmem_inst/mem_reg[11][0]  ( .D(n1025), .CK(clk), .Q(
        \xmem_inst/mem[11][0] ) );
  DFF_X1 \xmem_inst/mem_reg[11][1]  ( .D(n1024), .CK(clk), .Q(
        \xmem_inst/mem[11][1] ) );
  DFF_X1 \xmem_inst/mem_reg[11][2]  ( .D(n1023), .CK(clk), .Q(
        \xmem_inst/mem[11][2] ) );
  DFF_X1 \xmem_inst/mem_reg[11][3]  ( .D(n1022), .CK(clk), .Q(
        \xmem_inst/mem[11][3] ) );
  DFF_X1 \xmem_inst/mem_reg[11][4]  ( .D(n1021), .CK(clk), .Q(
        \xmem_inst/mem[11][4] ) );
  DFF_X1 \xmem_inst/mem_reg[11][5]  ( .D(n1020), .CK(clk), .Q(
        \xmem_inst/mem[11][5] ) );
  DFF_X1 \xmem_inst/mem_reg[11][6]  ( .D(n1019), .CK(clk), .Q(
        \xmem_inst/mem[11][6] ) );
  DFF_X1 \xmem_inst/mem_reg[11][7]  ( .D(n1018), .CK(clk), .Q(
        \xmem_inst/mem[11][7] ) );
  DFF_X1 \xmem_inst/mem_reg[11][8]  ( .D(n1017), .CK(clk), .Q(
        \xmem_inst/mem[11][8] ) );
  DFF_X1 \xmem_inst/mem_reg[11][9]  ( .D(n1016), .CK(clk), .Q(
        \xmem_inst/mem[11][9] ) );
  DFF_X1 \xmem_inst/mem_reg[11][10]  ( .D(n1015), .CK(clk), .Q(
        \xmem_inst/mem[11][10] ) );
  DFF_X1 \xmem_inst/mem_reg[12][0]  ( .D(n1014), .CK(clk), .Q(
        \xmem_inst/mem[12][0] ) );
  DFF_X1 \xmem_inst/mem_reg[12][1]  ( .D(n1013), .CK(clk), .Q(
        \xmem_inst/mem[12][1] ) );
  DFF_X1 \xmem_inst/mem_reg[12][2]  ( .D(n1012), .CK(clk), .Q(
        \xmem_inst/mem[12][2] ) );
  DFF_X1 \xmem_inst/mem_reg[12][3]  ( .D(n1011), .CK(clk), .Q(
        \xmem_inst/mem[12][3] ) );
  DFF_X1 \xmem_inst/mem_reg[12][4]  ( .D(n1010), .CK(clk), .Q(
        \xmem_inst/mem[12][4] ) );
  DFF_X1 \xmem_inst/mem_reg[12][5]  ( .D(n1009), .CK(clk), .Q(
        \xmem_inst/mem[12][5] ) );
  DFF_X1 \xmem_inst/mem_reg[12][6]  ( .D(n1008), .CK(clk), .Q(
        \xmem_inst/mem[12][6] ) );
  DFF_X1 \xmem_inst/mem_reg[12][7]  ( .D(n1007), .CK(clk), .Q(
        \xmem_inst/mem[12][7] ) );
  DFF_X1 \xmem_inst/mem_reg[12][8]  ( .D(n1006), .CK(clk), .Q(
        \xmem_inst/mem[12][8] ) );
  DFF_X1 \xmem_inst/mem_reg[12][9]  ( .D(n1005), .CK(clk), .Q(
        \xmem_inst/mem[12][9] ) );
  DFF_X1 \xmem_inst/mem_reg[12][10]  ( .D(n1004), .CK(clk), .Q(
        \xmem_inst/mem[12][10] ) );
  DFF_X1 \xmem_inst/mem_reg[13][0]  ( .D(n1003), .CK(clk), .Q(
        \xmem_inst/mem[13][0] ) );
  DFF_X1 \xmem_inst/mem_reg[13][1]  ( .D(n1002), .CK(clk), .Q(
        \xmem_inst/mem[13][1] ) );
  DFF_X1 \xmem_inst/mem_reg[13][2]  ( .D(n1001), .CK(clk), .Q(
        \xmem_inst/mem[13][2] ) );
  DFF_X1 \xmem_inst/mem_reg[13][3]  ( .D(n1000), .CK(clk), .Q(
        \xmem_inst/mem[13][3] ) );
  DFF_X1 \xmem_inst/mem_reg[13][4]  ( .D(n999), .CK(clk), .Q(
        \xmem_inst/mem[13][4] ) );
  DFF_X1 \xmem_inst/mem_reg[13][5]  ( .D(n998), .CK(clk), .Q(
        \xmem_inst/mem[13][5] ) );
  DFF_X1 \xmem_inst/mem_reg[13][6]  ( .D(n997), .CK(clk), .Q(
        \xmem_inst/mem[13][6] ) );
  DFF_X1 \xmem_inst/mem_reg[13][7]  ( .D(n996), .CK(clk), .Q(
        \xmem_inst/mem[13][7] ) );
  DFF_X1 \xmem_inst/mem_reg[13][8]  ( .D(n995), .CK(clk), .Q(
        \xmem_inst/mem[13][8] ) );
  DFF_X1 \xmem_inst/mem_reg[13][9]  ( .D(n994), .CK(clk), .Q(
        \xmem_inst/mem[13][9] ) );
  DFF_X1 \xmem_inst/mem_reg[13][10]  ( .D(n993), .CK(clk), .Q(
        \xmem_inst/mem[13][10] ) );
  DFF_X1 \xmem_inst/mem_reg[14][0]  ( .D(n992), .CK(clk), .Q(
        \xmem_inst/mem[14][0] ) );
  DFF_X1 \xmem_inst/mem_reg[14][1]  ( .D(n991), .CK(clk), .Q(
        \xmem_inst/mem[14][1] ) );
  DFF_X1 \xmem_inst/mem_reg[14][2]  ( .D(n990), .CK(clk), .Q(
        \xmem_inst/mem[14][2] ) );
  DFF_X1 \xmem_inst/mem_reg[14][3]  ( .D(n989), .CK(clk), .Q(
        \xmem_inst/mem[14][3] ) );
  DFF_X1 \xmem_inst/mem_reg[14][4]  ( .D(n988), .CK(clk), .Q(
        \xmem_inst/mem[14][4] ) );
  DFF_X1 \xmem_inst/mem_reg[14][5]  ( .D(n987), .CK(clk), .Q(
        \xmem_inst/mem[14][5] ) );
  DFF_X1 \xmem_inst/mem_reg[14][6]  ( .D(n986), .CK(clk), .Q(
        \xmem_inst/mem[14][6] ) );
  DFF_X1 \xmem_inst/mem_reg[14][7]  ( .D(n985), .CK(clk), .Q(
        \xmem_inst/mem[14][7] ) );
  DFF_X1 \xmem_inst/mem_reg[14][8]  ( .D(n984), .CK(clk), .Q(
        \xmem_inst/mem[14][8] ) );
  DFF_X1 \xmem_inst/mem_reg[14][9]  ( .D(n983), .CK(clk), .Q(
        \xmem_inst/mem[14][9] ) );
  DFF_X1 \xmem_inst/mem_reg[14][10]  ( .D(n982), .CK(clk), .Q(
        \xmem_inst/mem[14][10] ) );
  DFF_X1 \xmem_inst/mem_reg[15][0]  ( .D(n981), .CK(clk), .Q(
        \xmem_inst/mem[15][0] ) );
  DFF_X1 \xmem_inst/mem_reg[15][1]  ( .D(n980), .CK(clk), .Q(
        \xmem_inst/mem[15][1] ) );
  DFF_X1 \xmem_inst/mem_reg[15][2]  ( .D(n979), .CK(clk), .Q(
        \xmem_inst/mem[15][2] ) );
  DFF_X1 \xmem_inst/mem_reg[15][3]  ( .D(n978), .CK(clk), .Q(
        \xmem_inst/mem[15][3] ) );
  DFF_X1 \xmem_inst/mem_reg[15][4]  ( .D(n977), .CK(clk), .Q(
        \xmem_inst/mem[15][4] ) );
  DFF_X1 \xmem_inst/mem_reg[15][5]  ( .D(n976), .CK(clk), .Q(
        \xmem_inst/mem[15][5] ) );
  DFF_X1 \xmem_inst/mem_reg[15][6]  ( .D(n975), .CK(clk), .Q(
        \xmem_inst/mem[15][6] ) );
  DFF_X1 \xmem_inst/mem_reg[15][7]  ( .D(n974), .CK(clk), .Q(
        \xmem_inst/mem[15][7] ) );
  DFF_X1 \xmem_inst/mem_reg[15][8]  ( .D(n973), .CK(clk), .Q(
        \xmem_inst/mem[15][8] ) );
  DFF_X1 \xmem_inst/mem_reg[15][9]  ( .D(n972), .CK(clk), .Q(
        \xmem_inst/mem[15][9] ) );
  DFF_X1 \xmem_inst/mem_reg[15][10]  ( .D(n971), .CK(clk), .Q(
        \xmem_inst/mem[15][10] ) );
  DFF_X1 \xmem_inst/mem_reg[0][0]  ( .D(n1146), .CK(clk), .Q(
        \xmem_inst/mem[0][0] ) );
  DFF_X1 \xmem_inst/mem_reg[0][1]  ( .D(n1145), .CK(clk), .Q(
        \xmem_inst/mem[0][1] ) );
  DFF_X1 \xmem_inst/mem_reg[0][2]  ( .D(n1144), .CK(clk), .Q(
        \xmem_inst/mem[0][2] ) );
  DFF_X1 \xmem_inst/mem_reg[0][3]  ( .D(n1143), .CK(clk), .Q(
        \xmem_inst/mem[0][3] ) );
  DFF_X1 \xmem_inst/mem_reg[0][4]  ( .D(n1142), .CK(clk), .Q(
        \xmem_inst/mem[0][4] ) );
  DFF_X1 \xmem_inst/mem_reg[0][5]  ( .D(n1141), .CK(clk), .Q(
        \xmem_inst/mem[0][5] ) );
  DFF_X1 \xmem_inst/mem_reg[0][6]  ( .D(n1140), .CK(clk), .Q(
        \xmem_inst/mem[0][6] ) );
  DFF_X1 \xmem_inst/mem_reg[0][7]  ( .D(n1139), .CK(clk), .Q(
        \xmem_inst/mem[0][7] ) );
  DFF_X1 \xmem_inst/mem_reg[0][8]  ( .D(n1138), .CK(clk), .Q(
        \xmem_inst/mem[0][8] ) );
  DFF_X1 \xmem_inst/mem_reg[0][9]  ( .D(n1137), .CK(clk), .Q(
        \xmem_inst/mem[0][9] ) );
  DFF_X1 \xmem_inst/mem_reg[0][10]  ( .D(n1136), .CK(clk), .Q(
        \xmem_inst/mem[0][10] ) );
  DFF_X1 \xmem_inst/mem_reg[1][0]  ( .D(n1135), .CK(clk), .Q(
        \xmem_inst/mem[1][0] ) );
  DFF_X1 \xmem_inst/mem_reg[1][1]  ( .D(n1134), .CK(clk), .Q(
        \xmem_inst/mem[1][1] ) );
  DFF_X1 \xmem_inst/mem_reg[1][2]  ( .D(n1133), .CK(clk), .Q(
        \xmem_inst/mem[1][2] ) );
  DFF_X1 \xmem_inst/mem_reg[1][3]  ( .D(n1132), .CK(clk), .Q(
        \xmem_inst/mem[1][3] ) );
  DFF_X1 \xmem_inst/mem_reg[1][4]  ( .D(n1131), .CK(clk), .Q(
        \xmem_inst/mem[1][4] ) );
  DFF_X1 \xmem_inst/mem_reg[1][5]  ( .D(n1130), .CK(clk), .Q(
        \xmem_inst/mem[1][5] ) );
  DFF_X1 \xmem_inst/mem_reg[1][6]  ( .D(n1129), .CK(clk), .Q(
        \xmem_inst/mem[1][6] ) );
  DFF_X1 \xmem_inst/mem_reg[1][7]  ( .D(n1128), .CK(clk), .Q(
        \xmem_inst/mem[1][7] ) );
  DFF_X1 \xmem_inst/mem_reg[1][8]  ( .D(n1127), .CK(clk), .Q(
        \xmem_inst/mem[1][8] ) );
  DFF_X1 \xmem_inst/mem_reg[1][9]  ( .D(n1126), .CK(clk), .Q(
        \xmem_inst/mem[1][9] ) );
  DFF_X1 \xmem_inst/mem_reg[1][10]  ( .D(n1125), .CK(clk), .Q(
        \xmem_inst/mem[1][10] ) );
  DFF_X1 \xmem_inst/mem_reg[2][0]  ( .D(n1124), .CK(clk), .Q(
        \xmem_inst/mem[2][0] ) );
  DFF_X1 \xmem_inst/mem_reg[2][1]  ( .D(n1123), .CK(clk), .Q(
        \xmem_inst/mem[2][1] ) );
  DFF_X1 \xmem_inst/mem_reg[2][2]  ( .D(n1122), .CK(clk), .Q(
        \xmem_inst/mem[2][2] ) );
  DFF_X1 \xmem_inst/mem_reg[2][3]  ( .D(n1121), .CK(clk), .Q(
        \xmem_inst/mem[2][3] ) );
  DFF_X1 \xmem_inst/mem_reg[2][4]  ( .D(n1120), .CK(clk), .Q(
        \xmem_inst/mem[2][4] ) );
  DFF_X1 \xmem_inst/mem_reg[2][5]  ( .D(n1119), .CK(clk), .Q(
        \xmem_inst/mem[2][5] ) );
  DFF_X1 \xmem_inst/mem_reg[2][6]  ( .D(n1118), .CK(clk), .Q(
        \xmem_inst/mem[2][6] ) );
  DFF_X1 \xmem_inst/mem_reg[2][7]  ( .D(n1117), .CK(clk), .Q(
        \xmem_inst/mem[2][7] ) );
  DFF_X1 \xmem_inst/mem_reg[2][8]  ( .D(n1116), .CK(clk), .Q(
        \xmem_inst/mem[2][8] ) );
  DFF_X1 \xmem_inst/mem_reg[2][9]  ( .D(n1115), .CK(clk), .Q(
        \xmem_inst/mem[2][9] ) );
  DFF_X1 \xmem_inst/mem_reg[2][10]  ( .D(n1114), .CK(clk), .Q(
        \xmem_inst/mem[2][10] ) );
  DFF_X1 \xmem_inst/mem_reg[3][0]  ( .D(n1113), .CK(clk), .Q(
        \xmem_inst/mem[3][0] ) );
  DFF_X1 \xmem_inst/mem_reg[3][1]  ( .D(n1112), .CK(clk), .Q(
        \xmem_inst/mem[3][1] ) );
  DFF_X1 \xmem_inst/mem_reg[3][2]  ( .D(n1111), .CK(clk), .Q(
        \xmem_inst/mem[3][2] ) );
  DFF_X1 \xmem_inst/mem_reg[3][3]  ( .D(n1110), .CK(clk), .Q(
        \xmem_inst/mem[3][3] ) );
  DFF_X1 \xmem_inst/mem_reg[3][4]  ( .D(n1109), .CK(clk), .Q(
        \xmem_inst/mem[3][4] ) );
  DFF_X1 \xmem_inst/mem_reg[3][5]  ( .D(n1108), .CK(clk), .Q(
        \xmem_inst/mem[3][5] ) );
  DFF_X1 \xmem_inst/mem_reg[3][6]  ( .D(n1107), .CK(clk), .Q(
        \xmem_inst/mem[3][6] ) );
  DFF_X1 \xmem_inst/mem_reg[3][7]  ( .D(n1106), .CK(clk), .Q(
        \xmem_inst/mem[3][7] ) );
  DFF_X1 \xmem_inst/mem_reg[3][8]  ( .D(n1105), .CK(clk), .Q(
        \xmem_inst/mem[3][8] ) );
  DFF_X1 \xmem_inst/mem_reg[3][9]  ( .D(n1104), .CK(clk), .Q(
        \xmem_inst/mem[3][9] ) );
  DFF_X1 \xmem_inst/mem_reg[3][10]  ( .D(n1103), .CK(clk), .Q(
        \xmem_inst/mem[3][10] ) );
  DFF_X1 \xmem_inst/mem_reg[4][0]  ( .D(n1102), .CK(clk), .Q(
        \xmem_inst/mem[4][0] ) );
  DFF_X1 \xmem_inst/mem_reg[4][1]  ( .D(n1101), .CK(clk), .Q(
        \xmem_inst/mem[4][1] ) );
  DFF_X1 \xmem_inst/mem_reg[4][2]  ( .D(n1100), .CK(clk), .Q(
        \xmem_inst/mem[4][2] ) );
  DFF_X1 \xmem_inst/mem_reg[4][3]  ( .D(n1099), .CK(clk), .Q(
        \xmem_inst/mem[4][3] ) );
  DFF_X1 \xmem_inst/mem_reg[4][4]  ( .D(n1098), .CK(clk), .Q(
        \xmem_inst/mem[4][4] ) );
  DFF_X1 \xmem_inst/mem_reg[4][5]  ( .D(n1097), .CK(clk), .Q(
        \xmem_inst/mem[4][5] ) );
  DFF_X1 \xmem_inst/mem_reg[4][6]  ( .D(n1096), .CK(clk), .Q(
        \xmem_inst/mem[4][6] ) );
  DFF_X1 \xmem_inst/mem_reg[4][7]  ( .D(n1095), .CK(clk), .Q(
        \xmem_inst/mem[4][7] ) );
  DFF_X1 \xmem_inst/mem_reg[4][8]  ( .D(n1094), .CK(clk), .Q(
        \xmem_inst/mem[4][8] ) );
  DFF_X1 \xmem_inst/mem_reg[4][9]  ( .D(n1093), .CK(clk), .Q(
        \xmem_inst/mem[4][9] ) );
  DFF_X1 \xmem_inst/mem_reg[4][10]  ( .D(n1092), .CK(clk), .Q(
        \xmem_inst/mem[4][10] ) );
  DFF_X1 \xmem_inst/mem_reg[5][0]  ( .D(n1091), .CK(clk), .Q(
        \xmem_inst/mem[5][0] ) );
  DFF_X1 \xmem_inst/mem_reg[5][1]  ( .D(n1090), .CK(clk), .Q(
        \xmem_inst/mem[5][1] ) );
  DFF_X1 \xmem_inst/mem_reg[5][2]  ( .D(n1089), .CK(clk), .Q(
        \xmem_inst/mem[5][2] ) );
  DFF_X1 \xmem_inst/mem_reg[5][3]  ( .D(n1088), .CK(clk), .Q(
        \xmem_inst/mem[5][3] ) );
  DFF_X1 \xmem_inst/mem_reg[5][4]  ( .D(n1087), .CK(clk), .Q(
        \xmem_inst/mem[5][4] ) );
  DFF_X1 \xmem_inst/mem_reg[5][5]  ( .D(n1086), .CK(clk), .Q(
        \xmem_inst/mem[5][5] ) );
  DFF_X1 \xmem_inst/mem_reg[5][6]  ( .D(n1085), .CK(clk), .Q(
        \xmem_inst/mem[5][6] ) );
  DFF_X1 \xmem_inst/mem_reg[5][7]  ( .D(n1084), .CK(clk), .Q(
        \xmem_inst/mem[5][7] ) );
  DFF_X1 \xmem_inst/mem_reg[5][8]  ( .D(n1083), .CK(clk), .Q(
        \xmem_inst/mem[5][8] ) );
  DFF_X1 \xmem_inst/mem_reg[5][9]  ( .D(n1082), .CK(clk), .Q(
        \xmem_inst/mem[5][9] ) );
  DFF_X1 \xmem_inst/mem_reg[5][10]  ( .D(n1081), .CK(clk), .Q(
        \xmem_inst/mem[5][10] ) );
  DFF_X1 \xmem_inst/mem_reg[6][0]  ( .D(n1080), .CK(clk), .Q(
        \xmem_inst/mem[6][0] ) );
  DFF_X1 \xmem_inst/mem_reg[6][1]  ( .D(n1079), .CK(clk), .Q(
        \xmem_inst/mem[6][1] ) );
  DFF_X1 \xmem_inst/mem_reg[6][2]  ( .D(n1078), .CK(clk), .Q(
        \xmem_inst/mem[6][2] ) );
  DFF_X1 \xmem_inst/mem_reg[6][3]  ( .D(n1077), .CK(clk), .Q(
        \xmem_inst/mem[6][3] ) );
  DFF_X1 \xmem_inst/mem_reg[6][4]  ( .D(n1076), .CK(clk), .Q(
        \xmem_inst/mem[6][4] ) );
  DFF_X1 \xmem_inst/mem_reg[6][5]  ( .D(n1075), .CK(clk), .Q(
        \xmem_inst/mem[6][5] ) );
  DFF_X1 \xmem_inst/mem_reg[6][6]  ( .D(n1074), .CK(clk), .Q(
        \xmem_inst/mem[6][6] ) );
  DFF_X1 \xmem_inst/mem_reg[6][7]  ( .D(n1073), .CK(clk), .Q(
        \xmem_inst/mem[6][7] ) );
  DFF_X1 \xmem_inst/mem_reg[6][8]  ( .D(n1072), .CK(clk), .Q(
        \xmem_inst/mem[6][8] ) );
  DFF_X1 \xmem_inst/mem_reg[6][9]  ( .D(n1071), .CK(clk), .Q(
        \xmem_inst/mem[6][9] ) );
  DFF_X1 \xmem_inst/mem_reg[6][10]  ( .D(n1070), .CK(clk), .Q(
        \xmem_inst/mem[6][10] ) );
  DFF_X1 \xmem_inst/mem_reg[7][0]  ( .D(n1069), .CK(clk), .Q(
        \xmem_inst/mem[7][0] ) );
  DFF_X1 \xmem_inst/mem_reg[7][1]  ( .D(n1068), .CK(clk), .Q(
        \xmem_inst/mem[7][1] ) );
  DFF_X1 \xmem_inst/mem_reg[7][2]  ( .D(n1067), .CK(clk), .Q(
        \xmem_inst/mem[7][2] ) );
  DFF_X1 \xmem_inst/mem_reg[7][3]  ( .D(n1066), .CK(clk), .Q(
        \xmem_inst/mem[7][3] ) );
  DFF_X1 \xmem_inst/mem_reg[7][4]  ( .D(n1065), .CK(clk), .Q(
        \xmem_inst/mem[7][4] ) );
  DFF_X1 \xmem_inst/mem_reg[7][5]  ( .D(n1064), .CK(clk), .Q(
        \xmem_inst/mem[7][5] ) );
  DFF_X1 \xmem_inst/mem_reg[7][6]  ( .D(n1063), .CK(clk), .Q(
        \xmem_inst/mem[7][6] ) );
  DFF_X1 \xmem_inst/mem_reg[7][7]  ( .D(n1062), .CK(clk), .Q(
        \xmem_inst/mem[7][7] ) );
  DFF_X1 \xmem_inst/mem_reg[7][8]  ( .D(n1061), .CK(clk), .Q(
        \xmem_inst/mem[7][8] ) );
  DFF_X1 \xmem_inst/mem_reg[7][9]  ( .D(n1060), .CK(clk), .Q(
        \xmem_inst/mem[7][9] ) );
  DFF_X1 \xmem_inst/mem_reg[7][10]  ( .D(n1059), .CK(clk), .Q(
        \xmem_inst/mem[7][10] ) );
  DFF_X1 \xmem_inst/mem_reg[16][0]  ( .D(n970), .CK(clk), .Q(
        \xmem_inst/mem[16][0] ) );
  DFF_X1 \xmem_inst/mem_reg[16][1]  ( .D(n969), .CK(clk), .Q(
        \xmem_inst/mem[16][1] ) );
  DFF_X1 \xmem_inst/mem_reg[16][2]  ( .D(n968), .CK(clk), .Q(
        \xmem_inst/mem[16][2] ) );
  DFF_X1 \xmem_inst/mem_reg[16][3]  ( .D(n967), .CK(clk), .Q(
        \xmem_inst/mem[16][3] ) );
  DFF_X1 \xmem_inst/mem_reg[16][4]  ( .D(n966), .CK(clk), .Q(
        \xmem_inst/mem[16][4] ) );
  DFF_X1 \xmem_inst/mem_reg[16][5]  ( .D(n965), .CK(clk), .Q(
        \xmem_inst/mem[16][5] ) );
  DFF_X1 \xmem_inst/mem_reg[16][6]  ( .D(n964), .CK(clk), .Q(
        \xmem_inst/mem[16][6] ) );
  DFF_X1 \xmem_inst/mem_reg[16][7]  ( .D(n963), .CK(clk), .Q(
        \xmem_inst/mem[16][7] ) );
  DFF_X1 \xmem_inst/mem_reg[16][8]  ( .D(n962), .CK(clk), .Q(
        \xmem_inst/mem[16][8] ) );
  DFF_X1 \xmem_inst/mem_reg[16][9]  ( .D(n961), .CK(clk), .Q(
        \xmem_inst/mem[16][9] ) );
  DFF_X1 \xmem_inst/mem_reg[16][10]  ( .D(n960), .CK(clk), .Q(
        \xmem_inst/mem[16][10] ) );
  DFF_X1 \xmem_inst/mem_reg[17][0]  ( .D(n959), .CK(clk), .Q(
        \xmem_inst/mem[17][0] ) );
  DFF_X1 \xmem_inst/mem_reg[17][1]  ( .D(n958), .CK(clk), .Q(
        \xmem_inst/mem[17][1] ) );
  DFF_X1 \xmem_inst/mem_reg[17][2]  ( .D(n957), .CK(clk), .Q(
        \xmem_inst/mem[17][2] ) );
  DFF_X1 \xmem_inst/mem_reg[17][3]  ( .D(n956), .CK(clk), .Q(
        \xmem_inst/mem[17][3] ) );
  DFF_X1 \xmem_inst/mem_reg[17][4]  ( .D(n955), .CK(clk), .Q(
        \xmem_inst/mem[17][4] ) );
  DFF_X1 \xmem_inst/mem_reg[17][5]  ( .D(n954), .CK(clk), .Q(
        \xmem_inst/mem[17][5] ) );
  DFF_X1 \xmem_inst/mem_reg[17][6]  ( .D(n953), .CK(clk), .Q(
        \xmem_inst/mem[17][6] ) );
  DFF_X1 \xmem_inst/mem_reg[17][7]  ( .D(n952), .CK(clk), .Q(
        \xmem_inst/mem[17][7] ) );
  DFF_X1 \xmem_inst/mem_reg[17][8]  ( .D(n951), .CK(clk), .Q(
        \xmem_inst/mem[17][8] ) );
  DFF_X1 \xmem_inst/mem_reg[17][9]  ( .D(n950), .CK(clk), .Q(
        \xmem_inst/mem[17][9] ) );
  DFF_X1 \xmem_inst/mem_reg[17][10]  ( .D(n949), .CK(clk), .Q(
        \xmem_inst/mem[17][10] ) );
  DFF_X1 \xmem_inst/mem_reg[18][0]  ( .D(n948), .CK(clk), .Q(
        \xmem_inst/mem[18][0] ) );
  DFF_X1 \xmem_inst/mem_reg[18][1]  ( .D(n947), .CK(clk), .Q(
        \xmem_inst/mem[18][1] ) );
  DFF_X1 \xmem_inst/mem_reg[18][2]  ( .D(n946), .CK(clk), .Q(
        \xmem_inst/mem[18][2] ) );
  DFF_X1 \xmem_inst/mem_reg[18][3]  ( .D(n945), .CK(clk), .Q(
        \xmem_inst/mem[18][3] ) );
  DFF_X1 \xmem_inst/mem_reg[18][4]  ( .D(n944), .CK(clk), .Q(
        \xmem_inst/mem[18][4] ) );
  DFF_X1 \xmem_inst/mem_reg[18][5]  ( .D(n943), .CK(clk), .Q(
        \xmem_inst/mem[18][5] ) );
  DFF_X1 \xmem_inst/mem_reg[18][6]  ( .D(n942), .CK(clk), .Q(
        \xmem_inst/mem[18][6] ) );
  DFF_X1 \xmem_inst/mem_reg[18][7]  ( .D(n941), .CK(clk), .Q(
        \xmem_inst/mem[18][7] ) );
  DFF_X1 \xmem_inst/mem_reg[18][8]  ( .D(n940), .CK(clk), .Q(
        \xmem_inst/mem[18][8] ) );
  DFF_X1 \xmem_inst/mem_reg[18][9]  ( .D(n939), .CK(clk), .Q(
        \xmem_inst/mem[18][9] ) );
  DFF_X1 \xmem_inst/mem_reg[18][10]  ( .D(n938), .CK(clk), .Q(
        \xmem_inst/mem[18][10] ) );
  DFF_X1 \xmem_inst/mem_reg[19][0]  ( .D(n937), .CK(clk), .Q(
        \xmem_inst/mem[19][0] ) );
  DFF_X1 \xmem_inst/mem_reg[19][1]  ( .D(n936), .CK(clk), .Q(
        \xmem_inst/mem[19][1] ) );
  DFF_X1 \xmem_inst/mem_reg[19][2]  ( .D(n935), .CK(clk), .Q(
        \xmem_inst/mem[19][2] ) );
  DFF_X1 \xmem_inst/mem_reg[19][3]  ( .D(n934), .CK(clk), .Q(
        \xmem_inst/mem[19][3] ) );
  DFF_X1 \xmem_inst/mem_reg[19][4]  ( .D(n933), .CK(clk), .Q(
        \xmem_inst/mem[19][4] ) );
  DFF_X1 \xmem_inst/mem_reg[19][5]  ( .D(n932), .CK(clk), .Q(
        \xmem_inst/mem[19][5] ) );
  DFF_X1 \xmem_inst/mem_reg[19][6]  ( .D(n931), .CK(clk), .Q(
        \xmem_inst/mem[19][6] ) );
  DFF_X1 \xmem_inst/mem_reg[19][7]  ( .D(n930), .CK(clk), .Q(
        \xmem_inst/mem[19][7] ) );
  DFF_X1 \xmem_inst/mem_reg[19][8]  ( .D(n929), .CK(clk), .Q(
        \xmem_inst/mem[19][8] ) );
  DFF_X1 \xmem_inst/mem_reg[19][9]  ( .D(n928), .CK(clk), .Q(
        \xmem_inst/mem[19][9] ) );
  DFF_X1 \xmem_inst/mem_reg[19][10]  ( .D(n927), .CK(clk), .Q(
        \xmem_inst/mem[19][10] ) );
  DFF_X1 \xmem_inst/mem_reg[20][0]  ( .D(n926), .CK(clk), .Q(
        \xmem_inst/mem[20][0] ) );
  DFF_X1 \xmem_inst/mem_reg[20][1]  ( .D(n925), .CK(clk), .Q(
        \xmem_inst/mem[20][1] ) );
  DFF_X1 \xmem_inst/mem_reg[20][2]  ( .D(n924), .CK(clk), .Q(
        \xmem_inst/mem[20][2] ) );
  DFF_X1 \xmem_inst/mem_reg[20][3]  ( .D(n923), .CK(clk), .Q(
        \xmem_inst/mem[20][3] ) );
  DFF_X1 \xmem_inst/mem_reg[20][4]  ( .D(n922), .CK(clk), .Q(
        \xmem_inst/mem[20][4] ) );
  DFF_X1 \xmem_inst/mem_reg[20][5]  ( .D(n921), .CK(clk), .Q(
        \xmem_inst/mem[20][5] ) );
  DFF_X1 \xmem_inst/mem_reg[20][6]  ( .D(n920), .CK(clk), .Q(
        \xmem_inst/mem[20][6] ) );
  DFF_X1 \xmem_inst/mem_reg[20][7]  ( .D(n919), .CK(clk), .Q(
        \xmem_inst/mem[20][7] ) );
  DFF_X1 \xmem_inst/mem_reg[20][8]  ( .D(n918), .CK(clk), .Q(
        \xmem_inst/mem[20][8] ) );
  DFF_X1 \xmem_inst/mem_reg[20][9]  ( .D(n917), .CK(clk), .Q(
        \xmem_inst/mem[20][9] ) );
  DFF_X1 \xmem_inst/mem_reg[20][10]  ( .D(n916), .CK(clk), .Q(
        \xmem_inst/mem[20][10] ) );
  DFF_X1 \xmem_inst/mem_reg[21][0]  ( .D(n915), .CK(clk), .Q(
        \xmem_inst/mem[21][0] ) );
  DFF_X1 \xmem_inst/mem_reg[21][1]  ( .D(n914), .CK(clk), .Q(
        \xmem_inst/mem[21][1] ) );
  DFF_X1 \xmem_inst/mem_reg[21][2]  ( .D(n913), .CK(clk), .Q(
        \xmem_inst/mem[21][2] ) );
  DFF_X1 \xmem_inst/mem_reg[21][3]  ( .D(n912), .CK(clk), .Q(
        \xmem_inst/mem[21][3] ) );
  DFF_X1 \xmem_inst/mem_reg[21][4]  ( .D(n911), .CK(clk), .Q(
        \xmem_inst/mem[21][4] ) );
  DFF_X1 \xmem_inst/mem_reg[21][5]  ( .D(n910), .CK(clk), .Q(
        \xmem_inst/mem[21][5] ) );
  DFF_X1 \xmem_inst/mem_reg[21][6]  ( .D(n909), .CK(clk), .Q(
        \xmem_inst/mem[21][6] ) );
  DFF_X1 \xmem_inst/mem_reg[21][7]  ( .D(n908), .CK(clk), .Q(
        \xmem_inst/mem[21][7] ) );
  DFF_X1 \xmem_inst/mem_reg[21][8]  ( .D(n907), .CK(clk), .Q(
        \xmem_inst/mem[21][8] ) );
  DFF_X1 \xmem_inst/mem_reg[21][9]  ( .D(n906), .CK(clk), .Q(
        \xmem_inst/mem[21][9] ) );
  DFF_X1 \xmem_inst/mem_reg[21][10]  ( .D(n905), .CK(clk), .Q(
        \xmem_inst/mem[21][10] ) );
  DFF_X1 \xmem_inst/mem_reg[22][0]  ( .D(n904), .CK(clk), .Q(
        \xmem_inst/mem[22][0] ) );
  DFF_X1 \xmem_inst/mem_reg[22][1]  ( .D(n903), .CK(clk), .Q(
        \xmem_inst/mem[22][1] ) );
  DFF_X1 \xmem_inst/mem_reg[22][2]  ( .D(n902), .CK(clk), .Q(
        \xmem_inst/mem[22][2] ) );
  DFF_X1 \xmem_inst/mem_reg[22][3]  ( .D(n901), .CK(clk), .Q(
        \xmem_inst/mem[22][3] ) );
  DFF_X1 \xmem_inst/mem_reg[22][4]  ( .D(n900), .CK(clk), .Q(
        \xmem_inst/mem[22][4] ) );
  DFF_X1 \xmem_inst/mem_reg[22][5]  ( .D(n899), .CK(clk), .Q(
        \xmem_inst/mem[22][5] ) );
  DFF_X1 \xmem_inst/mem_reg[22][6]  ( .D(n898), .CK(clk), .Q(
        \xmem_inst/mem[22][6] ) );
  DFF_X1 \xmem_inst/mem_reg[22][7]  ( .D(n897), .CK(clk), .Q(
        \xmem_inst/mem[22][7] ) );
  DFF_X1 \xmem_inst/mem_reg[22][8]  ( .D(n896), .CK(clk), .Q(
        \xmem_inst/mem[22][8] ) );
  DFF_X1 \xmem_inst/mem_reg[22][9]  ( .D(n895), .CK(clk), .Q(
        \xmem_inst/mem[22][9] ) );
  DFF_X1 \xmem_inst/mem_reg[22][10]  ( .D(n894), .CK(clk), .Q(
        \xmem_inst/mem[22][10] ) );
  DFF_X1 \xmem_inst/mem_reg[23][0]  ( .D(n893), .CK(clk), .Q(
        \xmem_inst/mem[23][0] ) );
  DFF_X1 \xmem_inst/mem_reg[23][1]  ( .D(n892), .CK(clk), .Q(
        \xmem_inst/mem[23][1] ) );
  DFF_X1 \xmem_inst/mem_reg[23][2]  ( .D(n891), .CK(clk), .Q(
        \xmem_inst/mem[23][2] ) );
  DFF_X1 \xmem_inst/mem_reg[23][3]  ( .D(n890), .CK(clk), .Q(
        \xmem_inst/mem[23][3] ) );
  DFF_X1 \xmem_inst/mem_reg[23][4]  ( .D(n889), .CK(clk), .Q(
        \xmem_inst/mem[23][4] ) );
  DFF_X1 \xmem_inst/mem_reg[23][5]  ( .D(n888), .CK(clk), .Q(
        \xmem_inst/mem[23][5] ) );
  DFF_X1 \xmem_inst/mem_reg[23][6]  ( .D(n887), .CK(clk), .Q(
        \xmem_inst/mem[23][6] ) );
  DFF_X1 \xmem_inst/mem_reg[23][7]  ( .D(n886), .CK(clk), .Q(
        \xmem_inst/mem[23][7] ) );
  DFF_X1 \xmem_inst/mem_reg[23][8]  ( .D(n885), .CK(clk), .Q(
        \xmem_inst/mem[23][8] ) );
  DFF_X1 \xmem_inst/mem_reg[23][9]  ( .D(n884), .CK(clk), .Q(
        \xmem_inst/mem[23][9] ) );
  DFF_X1 \xmem_inst/mem_reg[23][10]  ( .D(n883), .CK(clk), .Q(
        \xmem_inst/mem[23][10] ) );
  DFF_X1 \fmem_addr_reg[0]  ( .D(n816), .CK(clk), .Q(fmem_addr[0]), .QN(n2496)
         );
  DFF_X1 \fmem_addr_reg[1]  ( .D(n815), .CK(clk), .Q(fmem_addr[1]), .QN(n2491)
         );
  DFF_X1 \fmem_addr_reg[2]  ( .D(n814), .CK(clk), .Q(fmem_addr[2]), .QN(n2489)
         );
  DFF_X1 \xmem_inst/mem_reg[29][0]  ( .D(n827), .CK(clk), .Q(
        \xmem_inst/mem[29][0] ) );
  DFF_X1 \xmem_inst/mem_reg[29][1]  ( .D(n826), .CK(clk), .Q(
        \xmem_inst/mem[29][1] ) );
  DFF_X1 \xmem_inst/mem_reg[29][2]  ( .D(n825), .CK(clk), .Q(
        \xmem_inst/mem[29][2] ) );
  DFF_X1 \xmem_inst/mem_reg[29][3]  ( .D(n824), .CK(clk), .Q(
        \xmem_inst/mem[29][3] ) );
  DFF_X1 \xmem_inst/mem_reg[29][4]  ( .D(n823), .CK(clk), .Q(
        \xmem_inst/mem[29][4] ) );
  DFF_X1 \xmem_inst/mem_reg[29][5]  ( .D(n822), .CK(clk), .Q(
        \xmem_inst/mem[29][5] ) );
  DFF_X1 \xmem_inst/mem_reg[29][6]  ( .D(n821), .CK(clk), .Q(
        \xmem_inst/mem[29][6] ) );
  DFF_X1 \xmem_inst/mem_reg[29][7]  ( .D(n820), .CK(clk), .Q(
        \xmem_inst/mem[29][7] ) );
  DFF_X1 \xmem_inst/mem_reg[29][8]  ( .D(n819), .CK(clk), .Q(
        \xmem_inst/mem[29][8] ) );
  DFF_X1 \xmem_inst/mem_reg[29][9]  ( .D(n818), .CK(clk), .Q(
        \xmem_inst/mem[29][9] ) );
  DFF_X1 \xmem_inst/mem_reg[29][10]  ( .D(n817), .CK(clk), .Q(
        \xmem_inst/mem[29][10] ) );
  DFF_X1 \ctrl_conv_output_inst/conv_start_accum_reg  ( .D(
        \ctrl_conv_output_inst/N74 ), .CK(clk), .QN(n2505) );
  DFF_X1 \fmem_inst/z_reg[1]  ( .D(n811), .CK(clk), .Q(fmem_data[1]), .QN(
        n2499) );
  DFF_X1 \fmem_inst/z_reg[4]  ( .D(n808), .CK(clk), .Q(fmem_data[4]), .QN(
        n2475) );
  DFF_X1 \fmem_inst/z_reg[3]  ( .D(n809), .CK(clk), .Q(fmem_data[3]), .QN(
        n2500) );
  DFF_X1 \fmem_inst/z_reg[10]  ( .D(n807), .CK(clk), .Q(fmem_data[10]), .QN(
        n2504) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[0]  ( .D(n794), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [0]), .QN(n2483) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[2]  ( .D(n792), .CK(clk), .Q(n2480) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[3]  ( .D(n791), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [3]) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[5]  ( .D(n789), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [5]) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[6]  ( .D(n788), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [6]) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[7]  ( .D(n787), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [7]), .QN(n1222) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[8]  ( .D(n786), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [8]) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[9]  ( .D(n785), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [9]) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[10]  ( .D(n784), .CK(clk), .QN(n2488) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[4]  ( .D(n801), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [4]), .QN(n2506) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[9]  ( .D(n796), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [9]), .QN(n2507) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[10]  ( .D(n795), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [10]), .QN(n2516) );
  DFF_X1 \fmem_addr_reg[3]  ( .D(n813), .CK(clk), .Q(fmem_addr[3]), .QN(n2498)
         );
  DFF_X1 \mac_unit_inst/adder_reg_reg[1]  ( .D(n793), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [1]), .QN(n2481) );
  DFF_X1 \mac_unit_inst/adder_reg_reg[4]  ( .D(n790), .CK(clk), .Q(
        \mac_unit_inst/adder_reg [4]) );
  DFF_X1 \xmem_inst/data_out_reg[10]  ( .D(\xmem_inst/N16 ), .CK(clk), .Q(
        xmem_data[10]), .QN(n2479) );
  DFF_X1 \xmem_inst/data_out_reg[3]  ( .D(n1233), .CK(clk), .Q(n2487), .QN(
        \DP_OP_65J1_122_2282/n664 ) );
  DFF_X1 \xmem_inst/data_out_reg[5]  ( .D(n1232), .CK(clk), .Q(n2478), .QN(
        \DP_OP_65J1_122_2282/n663 ) );
  DFF_X1 \xmem_inst/data_out_reg[9]  ( .D(n1220), .CK(clk), .Q(n2485), .QN(
        xmem_data[9]) );
  DFF_X1 \xmem_inst/data_out_reg[1]  ( .D(n1231), .CK(clk), .Q(n2473), .QN(
        xmem_data[1]) );
  DFF_X1 \xmem_inst/data_out_reg[0]  ( .D(n1230), .CK(clk), .Q(n2486), .QN(
        xmem_data[0]) );
  DFF_X1 \xmem_inst/data_out_reg[6]  ( .D(n1229), .CK(clk), .Q(n2484), .QN(
        xmem_data[6]) );
  DFF_X1 \ctrl_conv_output_inst/cnt_conv_reg[3]  ( .D(n2519), .CK(clk), .QN(
        \ctrl_conv_output_inst/cnt_conv [3]) );
  DFF_X1 \fmem_inst/z_reg[2]  ( .D(n2518), .CK(clk), .QN(fmem_data[2]) );
  SDFF_X1 \xmem_inst/data_out_reg[7]  ( .D(\xmem_inst/N19 ), .SI(1'b0), .SE(
        1'b0), .CK(clk), .Q(xmem_data[7]), .QN(n2476) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[1]  ( .D(n804), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [1]), .QN(n2517) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[2]  ( .D(n803), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [2]), .QN(n2508) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[0]  ( .D(n805), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [0]), .QN(n2520) );
  DFF_X1 \fmem_inst/z_reg[0]  ( .D(n812), .CK(clk), .Q(fmem_data[0]), .QN(
        n2494) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[6]  ( .D(n799), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [6]), .QN(n2509) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[7]  ( .D(n798), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [7]), .QN(n2510) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[8]  ( .D(n797), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [8]), .QN(n2513) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[3]  ( .D(n802), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [3]), .QN(n2514) );
  DFF_X1 \mac_unit_inst/x_mult_f_reg_reg[5]  ( .D(n800), .CK(clk), .Q(
        \mac_unit_inst/x_mult_f_reg [5]), .QN(n2515) );
  BUF_X1 U1187 ( .A(\DP_OP_65J1_122_2282/n663 ), .Z(n1205) );
  XOR2_X1 U1188 ( .A(n2473), .B(n2474), .Z(n1160) );
  AOI21_X1 U1189 ( .B1(n1512), .B2(n1913), .A(n1547), .ZN(n1750) );
  NAND2_X1 U1190 ( .A1(n2471), .A2(n2468), .ZN(n2465) );
  NOR2_X1 U1191 ( .A1(n2412), .A2(n2406), .ZN(n2467) );
  NOR2_X1 U1192 ( .A1(n1528), .A2(n1527), .ZN(n1340) );
  OR2_X1 U1193 ( .A1(n1464), .A2(n1171), .ZN(n1555) );
  OR2_X1 U1194 ( .A1(n1412), .A2(n1411), .ZN(n1175) );
  NOR2_X1 U1195 ( .A1(n1186), .A2(n1209), .ZN(n1509) );
  OAI21_X1 U1196 ( .B1(n1578), .B2(n1581), .A(n1579), .ZN(n1746) );
  OR2_X1 U1197 ( .A1(n1920), .A2(n2508), .ZN(n1576) );
  OR2_X1 U1198 ( .A1(n1920), .A2(n2514), .ZN(n1584) );
  OR2_X1 U1199 ( .A1(n1920), .A2(n2517), .ZN(n1569) );
  OR2_X1 U1200 ( .A1(n1279), .A2(n1278), .ZN(n1484) );
  OR2_X1 U1201 ( .A1(n1920), .A2(n2520), .ZN(n1562) );
  BUF_X1 U1202 ( .A(xmem_data[1]), .Z(n1395) );
  BUF_X1 U1203 ( .A(xmem_data[1]), .Z(n1372) );
  INV_X1 U1204 ( .A(n1529), .ZN(n1161) );
  AOI21_X1 U1205 ( .B1(n1467), .B2(n1466), .A(n1465), .ZN(n1162) );
  AOI21_X1 U1206 ( .B1(n1467), .B2(n1466), .A(n1465), .ZN(n1910) );
  INV_X1 U1207 ( .A(xmem_data[7]), .ZN(n1163) );
  BUF_X1 U1208 ( .A(n1915), .Z(n1164) );
  CLKBUF_X1 U1209 ( .A(n1294), .Z(n1194) );
  INV_X1 U1210 ( .A(n1191), .ZN(n1432) );
  INV_X1 U1211 ( .A(n1255), .ZN(n1249) );
  OR2_X1 U1212 ( .A1(n1324), .A2(n1269), .ZN(n1254) );
  NAND2_X1 U1213 ( .A1(n1371), .A2(fmem_data[0]), .ZN(n1384) );
  NAND2_X1 U1214 ( .A1(n1337), .A2(n1335), .ZN(n1308) );
  INV_X1 U1215 ( .A(n1310), .ZN(n1313) );
  CLKBUF_X1 U1216 ( .A(n1311), .Z(n1312) );
  NAND2_X1 U1217 ( .A1(n1366), .A2(n1365), .ZN(n1411) );
  AND2_X1 U1218 ( .A1(n2450), .A2(n1247), .ZN(n2401) );
  NAND2_X1 U1219 ( .A1(n1508), .A2(n1510), .ZN(n1913) );
  BUF_X1 U1220 ( .A(\DP_OP_65J1_122_2282/n664 ), .Z(n1203) );
  CLKBUF_X1 U1221 ( .A(n2478), .Z(n1165) );
  CLKBUF_X1 U1222 ( .A(\DP_OP_65J1_122_2282/n664 ), .Z(n1199) );
  NAND2_X1 U1223 ( .A1(n1302), .A2(n1301), .ZN(n1337) );
  INV_X1 U1224 ( .A(n1192), .ZN(n1299) );
  NAND2_X1 U1225 ( .A1(n1307), .A2(n1306), .ZN(n1335) );
  AND2_X1 U1226 ( .A1(n1272), .A2(fmem_data[0]), .ZN(n1310) );
  XNOR2_X1 U1227 ( .A(n1334), .B(n1333), .ZN(n1457) );
  NAND2_X1 U1228 ( .A1(n1319), .A2(n1318), .ZN(n1448) );
  OR2_X1 U1229 ( .A1(n1324), .A2(n1321), .ZN(n1318) );
  AND2_X1 U1230 ( .A1(fmem_data[0]), .A2(n1358), .ZN(n1413) );
  NAND3_X1 U1231 ( .A1(n1316), .A2(n1315), .A3(n1314), .ZN(n1518) );
  NAND2_X1 U1232 ( .A1(n1478), .A2(n1477), .ZN(n1504) );
  INV_X1 U1233 ( .A(n1474), .ZN(n1475) );
  CLKBUF_X1 U1234 ( .A(n1501), .Z(n1174) );
  INV_X1 U1235 ( .A(n1499), .ZN(n1500) );
  CLKBUF_X1 U1236 ( .A(n1420), .Z(n1204) );
  NAND2_X1 U1237 ( .A1(n1381), .A2(n1238), .ZN(n1409) );
  INV_X1 U1238 ( .A(n1384), .ZN(n1380) );
  XNOR2_X1 U1239 ( .A(n1347), .B(n1346), .ZN(n1521) );
  OR2_X1 U1240 ( .A1(n1507), .A2(n1506), .ZN(n1542) );
  CLKBUF_X1 U1241 ( .A(n1348), .Z(n1351) );
  NAND2_X1 U1242 ( .A1(n1454), .A2(n1453), .ZN(n1455) );
  INV_X1 U1243 ( .A(n1175), .ZN(n1550) );
  INV_X1 U1244 ( .A(n1172), .ZN(n1592) );
  INV_X1 U1245 ( .A(n1914), .ZN(n1512) );
  AOI21_X1 U1246 ( .B1(n2452), .B2(n2401), .A(n2400), .ZN(n2411) );
  INV_X1 U1247 ( .A(n2399), .ZN(n2400) );
  AOI21_X1 U1248 ( .B1(n2401), .B2(n2451), .A(n1245), .ZN(n2399) );
  INV_X1 U1249 ( .A(n2166), .ZN(n2276) );
  NAND2_X1 U1250 ( .A1(s_ready_x), .A2(s_valid_x), .ZN(n2166) );
  OR2_X1 U1251 ( .A1(n2166), .A2(n1938), .ZN(n2347) );
  INV_X1 U1252 ( .A(n1913), .ZN(n1749) );
  OR2_X1 U1253 ( .A1(n1750), .A2(n1225), .ZN(n1751) );
  NAND2_X1 U1254 ( .A1(n2381), .A2(n1944), .ZN(n1920) );
  NAND2_X1 U1255 ( .A1(n2456), .A2(\mac_unit_inst/adder_reg [8]), .ZN(n2459)
         );
  INV_X1 U1256 ( .A(n2475), .ZN(n1841) );
  INV_X1 U1257 ( .A(n2273), .ZN(n2272) );
  INV_X1 U1258 ( .A(n2069), .ZN(n2068) );
  INV_X1 U1259 ( .A(n2055), .ZN(n2054) );
  INV_X1 U1260 ( .A(n2163), .ZN(n2162) );
  AOI21_X1 U1261 ( .B1(n2464), .B2(n2454), .A(n1227), .ZN(n2455) );
  AND2_X1 U1262 ( .A1(n1911), .A2(n1246), .ZN(n1213) );
  AOI21_X1 U1263 ( .B1(n1201), .B2(n1491), .A(n1490), .ZN(n1166) );
  XNOR2_X1 U1264 ( .A(n1351), .B(n1167), .ZN(n1906) );
  XNOR2_X1 U1265 ( .A(n1350), .B(n1349), .ZN(n1167) );
  INV_X1 U1266 ( .A(n1197), .ZN(n1168) );
  AND2_X1 U1267 ( .A1(fmem_data[0]), .A2(n1501), .ZN(n1169) );
  AND2_X1 U1268 ( .A1(fmem_data[0]), .A2(n1501), .ZN(n1444) );
  NAND2_X1 U1269 ( .A1(n1258), .A2(n1257), .ZN(n1170) );
  XNOR2_X1 U1270 ( .A(n1460), .B(n1188), .ZN(n1171) );
  AND2_X1 U1271 ( .A1(n1412), .A2(n1411), .ZN(n1172) );
  XNOR2_X1 U1272 ( .A(n1289), .B(n1483), .ZN(n1173) );
  NAND2_X1 U1273 ( .A1(n1370), .A2(n1364), .ZN(n1366) );
  XNOR2_X1 U1274 ( .A(n1370), .B(n1369), .ZN(n1410) );
  OR2_X1 U1275 ( .A1(n1407), .A2(n1406), .ZN(n1745) );
  OAI21_X1 U1276 ( .B1(n1380), .B2(n1374), .A(n1383), .ZN(n1381) );
  XNOR2_X1 U1277 ( .A(xmem_data[7]), .B(n2484), .ZN(n1176) );
  XNOR2_X1 U1278 ( .A(n1345), .B(n1344), .ZN(n1347) );
  INV_X1 U1279 ( .A(n1468), .ZN(n1177) );
  AND2_X2 U1280 ( .A1(n1911), .A2(n1246), .ZN(n1178) );
  NAND2_X1 U1281 ( .A1(n1309), .A2(n1308), .ZN(n1350) );
  NAND2_X1 U1282 ( .A1(n1328), .A2(n1327), .ZN(n1179) );
  NAND2_X1 U1283 ( .A1(n1446), .A2(n1169), .ZN(n1180) );
  NAND2_X1 U1284 ( .A1(n1260), .A2(n1259), .ZN(n1181) );
  XNOR2_X1 U1285 ( .A(xmem_data[7]), .B(n2484), .ZN(n1425) );
  NAND2_X1 U1286 ( .A1(n1258), .A2(n1257), .ZN(n1290) );
  INV_X1 U1287 ( .A(n1211), .ZN(n1182) );
  INV_X1 U1288 ( .A(n1182), .ZN(n1183) );
  INV_X1 U1289 ( .A(n1182), .ZN(n1184) );
  INV_X1 U1290 ( .A(n1182), .ZN(n1185) );
  FA_X1 U1291 ( .A(n1497), .B(n1496), .CI(n1495), .S(n1186) );
  INV_X1 U1292 ( .A(n2504), .ZN(n1187) );
  BUF_X1 U1293 ( .A(n1459), .Z(n1188) );
  XNOR2_X1 U1294 ( .A(n2473), .B(n2474), .ZN(n1189) );
  XNOR2_X1 U1295 ( .A(n2473), .B(n2474), .ZN(n1190) );
  OR2_X1 U1296 ( .A1(n1415), .A2(n1414), .ZN(n1191) );
  XNOR2_X1 U1297 ( .A(n1368), .B(n1367), .ZN(n1369) );
  OR2_X1 U1298 ( .A1(n1368), .A2(n1367), .ZN(n1364) );
  NAND2_X1 U1299 ( .A1(n1368), .A2(n1367), .ZN(n1365) );
  XNOR2_X1 U1300 ( .A(xmem_data[7]), .B(n2500), .ZN(n1192) );
  OAI21_X1 U1301 ( .B1(n1502), .B2(n1174), .A(n1500), .ZN(n1503) );
  NAND2_X1 U1302 ( .A1(n1475), .A2(n1502), .ZN(n1478) );
  NAND2_X1 U1303 ( .A1(n1502), .A2(n1249), .ZN(n1252) );
  XNOR2_X1 U1304 ( .A(n2485), .B(n2499), .ZN(n1263) );
  NAND2_X1 U1305 ( .A1(n1294), .A2(n1295), .ZN(n1193) );
  NOR2_X1 U1306 ( .A1(n1464), .A2(n1463), .ZN(n1195) );
  NOR2_X1 U1307 ( .A1(n1464), .A2(n1463), .ZN(n1196) );
  XNOR2_X1 U1308 ( .A(n2487), .B(n2482), .ZN(n1211) );
  AND2_X1 U1309 ( .A1(n1274), .A2(n1273), .ZN(n1197) );
  BUF_X1 U1310 ( .A(n1325), .Z(n1198) );
  XOR2_X1 U1311 ( .A(n1554), .B(n1200), .Z(n1558) );
  AND2_X1 U1312 ( .A1(n1555), .A2(n1556), .ZN(n1200) );
  NOR2_X1 U1313 ( .A1(n1341), .A2(n1340), .ZN(n1201) );
  XNOR2_X1 U1314 ( .A(n1385), .B(n1384), .ZN(n1407) );
  OAI21_X2 U1315 ( .B1(n1915), .B2(n1749), .A(n1750), .ZN(n1561) );
  NAND2_X1 U1316 ( .A1(n1375), .A2(n1190), .ZN(n1202) );
  OR2_X1 U1317 ( .A1(n1420), .A2(n1419), .ZN(n1449) );
  OAI21_X1 U1318 ( .B1(n1207), .B2(n1586), .A(n1587), .ZN(n1206) );
  AOI21_X1 U1319 ( .B1(n1745), .B2(n1746), .A(n1408), .ZN(n1207) );
  AOI21_X1 U1320 ( .B1(n1745), .B2(n1746), .A(n1408), .ZN(n1208) );
  OAI21_X1 U1321 ( .B1(n1488), .B2(n1487), .A(n1486), .ZN(n1209) );
  XNOR2_X2 U1322 ( .A(n2476), .B(n2477), .ZN(n1250) );
  OAI21_X1 U1323 ( .B1(n1488), .B2(n1487), .A(n1486), .ZN(n1513) );
  INV_X1 U1324 ( .A(n1386), .ZN(n1210) );
  XNOR2_X1 U1325 ( .A(n2484), .B(n2478), .ZN(n1423) );
  NAND2_X1 U1326 ( .A1(n2456), .A2(\mac_unit_inst/x_mult_f_reg [8]), .ZN(n2458) );
  NOR2_X1 U1327 ( .A1(\mac_unit_inst/adder_reg [8]), .A2(
        \mac_unit_inst/x_mult_f_reg [8]), .ZN(n2397) );
  BUF_X1 U1328 ( .A(n1485), .Z(n1212) );
  XOR2_X1 U1329 ( .A(n1424), .B(n2494), .Z(n1323) );
  INV_X1 U1330 ( .A(n1180), .ZN(n1303) );
  AND2_X1 U1331 ( .A1(n1173), .A2(n1168), .ZN(n1530) );
  NOR2_X1 U1332 ( .A1(n1526), .A2(n1224), .ZN(n1214) );
  INV_X1 U1333 ( .A(n1169), .ZN(n1445) );
  OR2_X1 U1334 ( .A1(n1305), .A2(n1250), .ZN(n1306) );
  OR2_X1 U1335 ( .A1(n1250), .A2(n1499), .ZN(n1477) );
  NOR2_X1 U1336 ( .A1(n1516), .A2(n1532), .ZN(n1215) );
  OAI21_X1 U1337 ( .B1(n1217), .B2(n1749), .A(n1750), .ZN(n1216) );
  OAI21_X1 U1338 ( .B1(n1494), .B2(n1162), .A(n1166), .ZN(n1217) );
  XNOR2_X1 U1339 ( .A(n2478), .B(n1218), .ZN(n1294) );
  NOR2_X1 U1340 ( .A1(n1540), .A2(n1539), .ZN(n1219) );
  INV_X1 U1341 ( .A(n1547), .ZN(n1548) );
  NOR4_X1 U1342 ( .A1(n1703), .A2(n1702), .A3(n1701), .A4(n1700), .ZN(n1220)
         );
  XOR2_X1 U1343 ( .A(n1540), .B(n1539), .Z(n1221) );
  AND2_X1 U1344 ( .A1(\mac_unit_inst/x_mult_f_reg [7]), .A2(n2442), .ZN(n1223)
         );
  AND2_X1 U1345 ( .A1(n1518), .A2(n1905), .ZN(n1224) );
  XNOR2_X1 U1346 ( .A(xmem_data[9]), .B(n2479), .ZN(n1272) );
  NOR2_X1 U1347 ( .A1(n1920), .A2(n2506), .ZN(n1225) );
  OAI21_X1 U1348 ( .B1(n2452), .B2(n2451), .A(n2450), .ZN(n2456) );
  AND2_X1 U1349 ( .A1(n2462), .A2(\mac_unit_inst/adder_reg [3]), .ZN(n1226) );
  AND2_X1 U1350 ( .A1(n2462), .A2(\mac_unit_inst/adder_reg [8]), .ZN(n1227) );
  OR2_X1 U1351 ( .A1(n1454), .A2(n1453), .ZN(n1228) );
  NOR4_X1 U1352 ( .A1(n1643), .A2(n1642), .A3(n1641), .A4(n1640), .ZN(n1229)
         );
  NOR4_X1 U1353 ( .A1(n1663), .A2(n1662), .A3(n1661), .A4(n1660), .ZN(n1230)
         );
  NOR4_X1 U1354 ( .A1(n1683), .A2(n1682), .A3(n1681), .A4(n1680), .ZN(n1231)
         );
  NOR4_X1 U1355 ( .A1(n1723), .A2(n1722), .A3(n1721), .A4(n1720), .ZN(n1232)
         );
  NOR4_X1 U1356 ( .A1(n1743), .A2(n1742), .A3(n1741), .A4(n1740), .ZN(n1233)
         );
  XOR2_X1 U1357 ( .A(n1186), .B(n1209), .Z(n1234) );
  XOR2_X1 U1358 ( .A(n1543), .B(n1542), .Z(n1235) );
  OR2_X1 U1359 ( .A1(\mac_unit_inst/adder_reg [9]), .A2(
        \mac_unit_inst/x_mult_f_reg [9]), .ZN(n1236) );
  OR2_X1 U1360 ( .A1(\mac_unit_inst/adder_reg [4]), .A2(
        \mac_unit_inst/x_mult_f_reg [4]), .ZN(n1237) );
  OR2_X1 U1361 ( .A1(n1384), .A2(n1382), .ZN(n1238) );
  AND2_X1 U1362 ( .A1(n2462), .A2(\mac_unit_inst/adder_reg [9]), .ZN(n1239) );
  OR2_X1 U1363 ( .A1(n1920), .A2(n2515), .ZN(n1240) );
  OR2_X1 U1364 ( .A1(n1920), .A2(n2509), .ZN(n1241) );
  OR2_X1 U1365 ( .A1(n1920), .A2(n2510), .ZN(n1242) );
  OR2_X1 U1366 ( .A1(n1920), .A2(n2513), .ZN(n1243) );
  NAND2_X1 U1367 ( .A1(n1913), .A2(n1548), .ZN(n1244) );
  INV_X1 U1368 ( .A(n1250), .ZN(n1501) );
  NAND2_X1 U1369 ( .A1(n1236), .A2(n2398), .ZN(n1245) );
  AND2_X1 U1370 ( .A1(n1912), .A2(n1548), .ZN(n1246) );
  AND2_X1 U1371 ( .A1(n2396), .A2(n2457), .ZN(n1247) );
  OR2_X1 U1372 ( .A1(n1749), .A2(n1225), .ZN(n1248) );
  XNOR2_X1 U1374 ( .A(n2477), .B(xmem_data[9]), .ZN(n1304) );
  AND2_X2 U1375 ( .A1(n1250), .A2(n1304), .ZN(n1502) );
  XNOR2_X1 U1376 ( .A(xmem_data[9]), .B(fmem_data[2]), .ZN(n1255) );
  XNOR2_X1 U1377 ( .A(xmem_data[9]), .B(fmem_data[3]), .ZN(n1284) );
  OR2_X1 U1378 ( .A1(n1250), .A2(n1284), .ZN(n1251) );
  NAND2_X1 U1379 ( .A1(n1252), .A2(n1251), .ZN(n1279) );
  XNOR2_X1 U1380 ( .A(\DP_OP_65J1_122_2282/n663 ), .B(xmem_data[6]), .ZN(n1421) );
  NAND2_X1 U1381 ( .A1(n1176), .A2(n1421), .ZN(n1324) );
  XNOR2_X1 U1382 ( .A(xmem_data[7]), .B(fmem_data[4]), .ZN(n1269) );
  XNOR2_X1 U1383 ( .A(n1424), .B(fmem_data[10]), .ZN(n1281) );
  OR2_X1 U1384 ( .A1(n1421), .A2(n1281), .ZN(n1253) );
  NAND2_X1 U1385 ( .A1(n1254), .A2(n1253), .ZN(n1278) );
  XNOR2_X1 U1386 ( .A(n1279), .B(n1278), .ZN(n1344) );
  OR2_X1 U1387 ( .A1(n1250), .A2(n1255), .ZN(n1258) );
  INV_X1 U1388 ( .A(n1263), .ZN(n1256) );
  NAND3_X1 U1389 ( .A1(n1304), .A2(n1256), .A3(n1250), .ZN(n1257) );
  XNOR2_X1 U1390 ( .A(n2487), .B(n2482), .ZN(n1295) );
  NAND2_X1 U1391 ( .A1(n1294), .A2(n1295), .ZN(n1429) );
  NAND2_X1 U1392 ( .A1(n1429), .A2(n1183), .ZN(n1260) );
  XNOR2_X1 U1393 ( .A(n1205), .B(fmem_data[10]), .ZN(n1261) );
  INV_X1 U1394 ( .A(n1261), .ZN(n1259) );
  NAND2_X1 U1395 ( .A1(n1260), .A2(n1259), .ZN(n1291) );
  OR2_X1 U1396 ( .A1(n1185), .A2(n1261), .ZN(n1332) );
  INV_X1 U1397 ( .A(n2485), .ZN(n1476) );
  XOR2_X1 U1398 ( .A(n1476), .B(fmem_data[0]), .Z(n1262) );
  NAND2_X1 U1399 ( .A1(n1262), .A2(n1502), .ZN(n1330) );
  OR2_X1 U1400 ( .A1(n1250), .A2(n1263), .ZN(n1329) );
  XNOR2_X1 U1401 ( .A(\DP_OP_65J1_122_2282/n663 ), .B(fmem_data[4]), .ZN(n1296) );
  INV_X1 U1402 ( .A(n1296), .ZN(n1264) );
  NAND3_X1 U1403 ( .A1(n1185), .A2(n1194), .A3(n1264), .ZN(n1331) );
  NAND4_X1 U1404 ( .A1(n1332), .A2(n1330), .A3(n1329), .A4(n1331), .ZN(n1292)
         );
  OAI21_X1 U1405 ( .B1(n1170), .B2(n1181), .A(n1292), .ZN(n1266) );
  NAND2_X1 U1406 ( .A1(n1181), .A2(n1170), .ZN(n1265) );
  NAND2_X1 U1407 ( .A1(n1266), .A2(n1265), .ZN(n1345) );
  OR2_X1 U1408 ( .A1(fmem_data[0]), .A2(n2479), .ZN(n1267) );
  INV_X1 U1409 ( .A(n1272), .ZN(n1506) );
  NOR2_X1 U1410 ( .A1(n1267), .A2(n1506), .ZN(n1277) );
  XNOR2_X1 U1411 ( .A(xmem_data[10]), .B(fmem_data[1]), .ZN(n1268) );
  NOR2_X1 U1412 ( .A1(n1268), .A2(n1506), .ZN(n1276) );
  NAND3_X1 U1413 ( .A1(n1192), .A2(n1423), .A3(n1425), .ZN(n1271) );
  XNOR2_X1 U1414 ( .A(\DP_OP_65J1_122_2282/n663 ), .B(xmem_data[6]), .ZN(n1280) );
  OR2_X1 U1415 ( .A1(n1269), .A2(n1280), .ZN(n1270) );
  NAND2_X1 U1416 ( .A1(n1271), .A2(n1270), .ZN(n1311) );
  AND2_X1 U1417 ( .A1(n1311), .A2(n1310), .ZN(n1275) );
  OAI21_X1 U1418 ( .B1(n1344), .B2(n1345), .A(n1346), .ZN(n1274) );
  NAND2_X1 U1419 ( .A1(n1345), .A2(n1344), .ZN(n1273) );
  NAND2_X1 U1420 ( .A1(n1274), .A2(n1273), .ZN(n1527) );
  FA_X1 U1421 ( .A(n1277), .B(n1276), .CI(n1275), .CO(n1485), .S(n1346) );
  XNOR2_X1 U1422 ( .A(n1485), .B(n1484), .ZN(n1289) );
  INV_X1 U1423 ( .A(n1280), .ZN(n1358) );
  OR2_X1 U1424 ( .A1(n1425), .A2(n1358), .ZN(n1283) );
  INV_X1 U1425 ( .A(n1281), .ZN(n1282) );
  NAND2_X1 U1426 ( .A1(n1282), .A2(n1283), .ZN(n1482) );
  INV_X1 U1427 ( .A(n1284), .ZN(n1285) );
  NAND3_X1 U1428 ( .A1(n1285), .A2(n1250), .A3(n1304), .ZN(n1287) );
  XNOR2_X1 U1429 ( .A(xmem_data[9]), .B(n1841), .ZN(n1474) );
  OR2_X1 U1430 ( .A1(n1474), .A2(n1250), .ZN(n1286) );
  NAND2_X1 U1431 ( .A1(n1287), .A2(n1286), .ZN(n1481) );
  XNOR2_X1 U1432 ( .A(xmem_data[10]), .B(fmem_data[2]), .ZN(n1288) );
  NOR2_X1 U1433 ( .A1(n1288), .A2(n1506), .ZN(n1480) );
  XNOR2_X1 U1434 ( .A(n1289), .B(n1483), .ZN(n1528) );
  XNOR2_X1 U1435 ( .A(n1527), .B(n1173), .ZN(n1473) );
  XNOR2_X1 U1436 ( .A(n1291), .B(n1290), .ZN(n1293) );
  XNOR2_X1 U1437 ( .A(n1293), .B(n1292), .ZN(n1348) );
  XNOR2_X1 U1438 ( .A(\DP_OP_65J1_122_2282/n663 ), .B(n2500), .ZN(n1428) );
  NAND3_X1 U1439 ( .A1(n1294), .A2(n1428), .A3(n1295), .ZN(n1298) );
  OR2_X1 U1440 ( .A1(n1296), .A2(n1211), .ZN(n1297) );
  NAND2_X1 U1441 ( .A1(n1298), .A2(n1297), .ZN(n1446) );
  NAND2_X1 U1442 ( .A1(n1446), .A2(n1444), .ZN(n1336) );
  OR2_X1 U1443 ( .A1(n1299), .A2(n1421), .ZN(n1302) );
  XNOR2_X1 U1444 ( .A(n1424), .B(fmem_data[2]), .ZN(n1317) );
  INV_X1 U1445 ( .A(n1317), .ZN(n1300) );
  NAND3_X1 U1446 ( .A1(n1425), .A2(n1300), .A3(n1423), .ZN(n1301) );
  NAND2_X1 U1447 ( .A1(n1303), .A2(n1337), .ZN(n1309) );
  NAND3_X1 U1448 ( .A1(n1304), .A2(n1250), .A3(n1476), .ZN(n1307) );
  OR2_X1 U1449 ( .A1(fmem_data[0]), .A2(n2485), .ZN(n1305) );
  NAND2_X1 U1450 ( .A1(n1348), .A2(n1350), .ZN(n1316) );
  XNOR2_X1 U1451 ( .A(n1313), .B(n1312), .ZN(n1349) );
  NAND2_X1 U1452 ( .A1(n1348), .A2(n1349), .ZN(n1315) );
  NAND2_X1 U1453 ( .A1(n1350), .A2(n1349), .ZN(n1314) );
  OR2_X1 U1454 ( .A1(n1423), .A2(n1317), .ZN(n1319) );
  XNOR2_X1 U1455 ( .A(xmem_data[7]), .B(fmem_data[1]), .ZN(n1321) );
  INV_X1 U1456 ( .A(n1160), .ZN(n1392) );
  XOR2_X1 U1457 ( .A(\DP_OP_65J1_122_2282/n664 ), .B(xmem_data[2]), .Z(n1375)
         );
  NAND2_X1 U1458 ( .A1(n1375), .A2(n1190), .ZN(n1394) );
  XNOR2_X1 U1459 ( .A(fmem_data[10]), .B(n1203), .ZN(n1325) );
  AOI21_X1 U1460 ( .B1(n1392), .B2(n1394), .A(n1198), .ZN(n1320) );
  INV_X1 U1461 ( .A(n1320), .ZN(n1447) );
  OR2_X1 U1462 ( .A1(n1423), .A2(n1321), .ZN(n1322) );
  OAI21_X1 U1463 ( .B1(n1324), .B2(n1323), .A(n1322), .ZN(n1420) );
  XNOR2_X1 U1464 ( .A(n1203), .B(n1841), .ZN(n1356) );
  OR2_X1 U1465 ( .A1(n1325), .A2(n1189), .ZN(n1326) );
  OAI21_X1 U1466 ( .B1(n1394), .B2(n1356), .A(n1326), .ZN(n1419) );
  OAI21_X1 U1467 ( .B1(n1448), .B2(n1447), .A(n1449), .ZN(n1328) );
  NAND2_X1 U1468 ( .A1(n1447), .A2(n1448), .ZN(n1327) );
  NAND2_X1 U1469 ( .A1(n1328), .A2(n1327), .ZN(n1458) );
  NAND2_X1 U1470 ( .A1(n1330), .A2(n1329), .ZN(n1334) );
  NAND2_X1 U1471 ( .A1(n1332), .A2(n1331), .ZN(n1333) );
  XNOR2_X1 U1472 ( .A(n1336), .B(n1335), .ZN(n1339) );
  INV_X1 U1473 ( .A(n1337), .ZN(n1338) );
  XNOR2_X1 U1474 ( .A(n1339), .B(n1338), .ZN(n1459) );
  OAI21_X1 U1475 ( .B1(n1458), .B2(n1457), .A(n1459), .ZN(n1343) );
  NAND2_X1 U1476 ( .A1(n1179), .A2(n1457), .ZN(n1342) );
  NAND2_X1 U1477 ( .A1(n1343), .A2(n1342), .ZN(n1905) );
  OR2_X1 U1478 ( .A1(n1518), .A2(n1905), .ZN(n1472) );
  NOR2_X1 U1479 ( .A1(n1473), .A2(n1472), .ZN(n1341) );
  NOR2_X1 U1480 ( .A1(n1341), .A2(n1340), .ZN(n1492) );
  NAND2_X1 U1481 ( .A1(n1343), .A2(n1342), .ZN(n1517) );
  XNOR2_X1 U1482 ( .A(n1518), .B(n1517), .ZN(n1469) );
  NOR2_X1 U1483 ( .A1(n1469), .A2(n1521), .ZN(n1471) );
  INV_X1 U1484 ( .A(n1905), .ZN(n1468) );
  NOR2_X1 U1485 ( .A1(n1906), .A2(n1468), .ZN(n1519) );
  NOR2_X1 U1486 ( .A1(n1471), .A2(n1519), .ZN(n1352) );
  NAND2_X1 U1487 ( .A1(n1492), .A2(n1352), .ZN(n1494) );
  OR2_X1 U1488 ( .A1(fmem_data[0]), .A2(n1165), .ZN(n1353) );
  OAI22_X1 U1489 ( .A1(n1193), .A2(n1165), .B1(n1353), .B2(n1184), .ZN(n1362)
         );
  XNOR2_X1 U1490 ( .A(n1205), .B(fmem_data[0]), .ZN(n1354) );
  XNOR2_X1 U1491 ( .A(n1205), .B(fmem_data[1]), .ZN(n1355) );
  OAI22_X1 U1492 ( .A1(n1193), .A2(n1354), .B1(n1184), .B2(n1355), .ZN(n1361)
         );
  XNOR2_X1 U1493 ( .A(n1205), .B(fmem_data[2]), .ZN(n1430) );
  OAI22_X1 U1494 ( .A1(n1193), .A2(n1355), .B1(n1184), .B2(n1430), .ZN(n1434)
         );
  INV_X1 U1495 ( .A(n2487), .ZN(n1386) );
  XNOR2_X1 U1496 ( .A(n1386), .B(fmem_data[3]), .ZN(n1363) );
  OR2_X1 U1497 ( .A1(n1190), .A2(n1356), .ZN(n1357) );
  OAI21_X1 U1498 ( .B1(n1394), .B2(n1363), .A(n1357), .ZN(n1416) );
  XNOR2_X1 U1499 ( .A(n1187), .B(n1372), .ZN(n1415) );
  INV_X1 U1500 ( .A(n1372), .ZN(n1397) );
  AND2_X1 U1501 ( .A1(n1397), .A2(n2486), .ZN(n1414) );
  NOR2_X1 U1502 ( .A1(n1415), .A2(n1414), .ZN(n1359) );
  XNOR2_X1 U1503 ( .A(n1413), .B(n1359), .ZN(n1360) );
  XNOR2_X1 U1504 ( .A(n1360), .B(n1416), .ZN(n1433) );
  HA_X1 U1505 ( .A(n1362), .B(n1361), .CO(n1435), .S(n1370) );
  XNOR2_X1 U1506 ( .A(n1199), .B(fmem_data[2]), .ZN(n1377) );
  OAI22_X1 U1507 ( .A1(n1202), .A2(n1377), .B1(n1363), .B2(n1392), .ZN(n1368)
         );
  NAND2_X1 U1508 ( .A1(n2486), .A2(n1395), .ZN(n1400) );
  XNOR2_X1 U1509 ( .A(n1372), .B(n1841), .ZN(n1373) );
  OAI22_X1 U1510 ( .A1(n1400), .A2(n1373), .B1(n1415), .B2(n2486), .ZN(n1367)
         );
  INV_X1 U1511 ( .A(n1185), .ZN(n1371) );
  XNOR2_X1 U1512 ( .A(n1395), .B(fmem_data[3]), .ZN(n1389) );
  OAI22_X1 U1513 ( .A1(n1400), .A2(n1389), .B1(n1373), .B2(n2486), .ZN(n1374)
         );
  INV_X1 U1514 ( .A(n1374), .ZN(n1382) );
  XNOR2_X1 U1515 ( .A(n1199), .B(fmem_data[1]), .ZN(n1387) );
  INV_X1 U1516 ( .A(n1387), .ZN(n1376) );
  NAND3_X1 U1517 ( .A1(n1376), .A2(n1375), .A3(n1189), .ZN(n1379) );
  OR2_X1 U1518 ( .A1(n1377), .A2(n1189), .ZN(n1378) );
  NAND2_X1 U1519 ( .A1(n1379), .A2(n1378), .ZN(n1383) );
  NOR2_X1 U1520 ( .A1(n1410), .A2(n1409), .ZN(n1586) );
  XNOR2_X1 U1521 ( .A(n1383), .B(n1382), .ZN(n1385) );
  XNOR2_X1 U1522 ( .A(n1386), .B(fmem_data[0]), .ZN(n1388) );
  OAI22_X1 U1523 ( .A1(n1202), .A2(n1388), .B1(n1387), .B2(n1392), .ZN(n1391)
         );
  XNOR2_X1 U1524 ( .A(n1395), .B(fmem_data[2]), .ZN(n1396) );
  OAI22_X1 U1525 ( .A1(n1400), .A2(n1396), .B1(n1389), .B2(n2486), .ZN(n1390)
         );
  HA_X1 U1526 ( .A(n1391), .B(n1390), .CO(n1406), .S(n1405) );
  OR2_X1 U1527 ( .A1(fmem_data[0]), .A2(n1210), .ZN(n1393) );
  OAI22_X1 U1528 ( .A1(n1202), .A2(n1210), .B1(n1393), .B2(n1392), .ZN(n1404)
         );
  NOR2_X1 U1529 ( .A1(n1405), .A2(n1404), .ZN(n1578) );
  XNOR2_X1 U1530 ( .A(n1395), .B(fmem_data[1]), .ZN(n1399) );
  OAI22_X1 U1531 ( .A1(n1400), .A2(n1399), .B1(n1396), .B2(n2486), .ZN(n1402)
         );
  AND2_X1 U1532 ( .A1(fmem_data[0]), .A2(n1160), .ZN(n1401) );
  OR2_X1 U1533 ( .A1(n1402), .A2(n1401), .ZN(n1572) );
  OR2_X1 U1534 ( .A1(fmem_data[0]), .A2(n1397), .ZN(n1398) );
  NAND2_X1 U1535 ( .A1(n1398), .A2(n1400), .ZN(n1565) );
  OAI22_X1 U1536 ( .A1(n1400), .A2(fmem_data[0]), .B1(n1399), .B2(n2486), .ZN(
        n1564) );
  NAND2_X1 U1537 ( .A1(n1565), .A2(n1564), .ZN(n1566) );
  INV_X1 U1538 ( .A(n1566), .ZN(n1573) );
  NAND2_X1 U1539 ( .A1(n1402), .A2(n1401), .ZN(n1571) );
  INV_X1 U1540 ( .A(n1571), .ZN(n1403) );
  AOI21_X1 U1541 ( .B1(n1572), .B2(n1573), .A(n1403), .ZN(n1581) );
  NAND2_X1 U1542 ( .A1(n1405), .A2(n1404), .ZN(n1579) );
  NAND2_X1 U1543 ( .A1(n1407), .A2(n1406), .ZN(n1744) );
  INV_X1 U1544 ( .A(n1744), .ZN(n1408) );
  NAND2_X1 U1545 ( .A1(n1410), .A2(n1409), .ZN(n1587) );
  OAI21_X1 U1546 ( .B1(n1586), .B2(n1208), .A(n1587), .ZN(n1549) );
  AOI21_X1 U1547 ( .B1(n1206), .B2(n1175), .A(n1172), .ZN(n1438) );
  OAI21_X1 U1548 ( .B1(n1413), .B2(n1432), .A(n1416), .ZN(n1418) );
  NAND2_X1 U1549 ( .A1(n1413), .A2(n1432), .ZN(n1417) );
  NAND2_X1 U1550 ( .A1(n1418), .A2(n1417), .ZN(n1441) );
  XNOR2_X1 U1551 ( .A(n1204), .B(n1419), .ZN(n1440) );
  OR2_X1 U1552 ( .A1(fmem_data[0]), .A2(n1163), .ZN(n1422) );
  OR2_X1 U1553 ( .A1(n1421), .A2(n1422), .ZN(n1427) );
  INV_X1 U1554 ( .A(n2476), .ZN(n1424) );
  NAND3_X1 U1555 ( .A1(n1176), .A2(n1424), .A3(n1423), .ZN(n1426) );
  NAND2_X1 U1556 ( .A1(n1427), .A2(n1426), .ZN(n1443) );
  INV_X1 U1557 ( .A(n1428), .ZN(n1431) );
  OAI22_X1 U1558 ( .A1(n1184), .A2(n1431), .B1(n1429), .B2(n1430), .ZN(n1442)
         );
  FA_X1 U1559 ( .A(n1435), .B(n1434), .CI(n1433), .CO(n1436), .S(n1412) );
  NOR2_X1 U1560 ( .A1(n1437), .A2(n1436), .ZN(n1597) );
  NAND2_X1 U1561 ( .A1(n1437), .A2(n1436), .ZN(n1603) );
  OAI21_X1 U1562 ( .B1(n1438), .B2(n1597), .A(n1603), .ZN(n1467) );
  FA_X1 U1563 ( .A(n1441), .B(n1440), .CI(n1439), .CO(n1461), .S(n1437) );
  FA_X1 U1564 ( .A(n1191), .B(n1443), .CI(n1442), .CO(n1454), .S(n1439) );
  XNOR2_X1 U1565 ( .A(n1446), .B(n1445), .ZN(n1453) );
  XNOR2_X1 U1566 ( .A(n1454), .B(n1453), .ZN(n1451) );
  XNOR2_X1 U1567 ( .A(n1448), .B(n1447), .ZN(n1450) );
  XNOR2_X1 U1568 ( .A(n1450), .B(n1449), .ZN(n1452) );
  XNOR2_X1 U1569 ( .A(n1452), .B(n1451), .ZN(n1462) );
  NOR2_X1 U1570 ( .A1(n1461), .A2(n1462), .ZN(n1607) );
  NAND2_X1 U1571 ( .A1(n1228), .A2(n1452), .ZN(n1456) );
  NAND2_X1 U1572 ( .A1(n1456), .A2(n1455), .ZN(n1464) );
  XNOR2_X1 U1573 ( .A(n1179), .B(n1457), .ZN(n1460) );
  XNOR2_X1 U1574 ( .A(n1460), .B(n1188), .ZN(n1463) );
  NOR2_X1 U1575 ( .A1(n1195), .A2(n1607), .ZN(n1466) );
  NAND2_X1 U1576 ( .A1(n1462), .A2(n1461), .ZN(n1608) );
  NAND2_X1 U1577 ( .A1(n1464), .A2(n1171), .ZN(n1556) );
  OAI21_X1 U1578 ( .B1(n1196), .B2(n1608), .A(n1556), .ZN(n1465) );
  NAND2_X1 U1579 ( .A1(n1906), .A2(n1468), .ZN(n1524) );
  NAND2_X1 U1580 ( .A1(n1469), .A2(n1521), .ZN(n1470) );
  OAI21_X1 U1581 ( .B1(n1471), .B2(n1524), .A(n1470), .ZN(n1491) );
  NAND2_X1 U1582 ( .A1(n1473), .A2(n1472), .ZN(n1489) );
  XNOR2_X1 U1583 ( .A(fmem_data[10]), .B(n1476), .ZN(n1499) );
  INV_X1 U1584 ( .A(n1504), .ZN(n1497) );
  XNOR2_X1 U1585 ( .A(xmem_data[10]), .B(fmem_data[3]), .ZN(n1479) );
  NOR2_X1 U1586 ( .A1(n1479), .A2(n1506), .ZN(n1496) );
  FA_X1 U1587 ( .A(n1482), .B(n1480), .CI(n1481), .CO(n1495), .S(n1483) );
  INV_X1 U1588 ( .A(n1483), .ZN(n1488) );
  NOR2_X1 U1589 ( .A1(n1212), .A2(n1484), .ZN(n1487) );
  NAND2_X1 U1590 ( .A1(n1212), .A2(n1484), .ZN(n1486) );
  OAI21_X1 U1591 ( .B1(n1340), .B2(n1489), .A(n1234), .ZN(n1490) );
  AOI21_X1 U1592 ( .B1(n1201), .B2(n1491), .A(n1490), .ZN(n1493) );
  OAI21_X1 U1593 ( .B1(n1494), .B2(n1910), .A(n1493), .ZN(n1915) );
  FA_X1 U1594 ( .A(n1497), .B(n1496), .CI(n1495), .CO(n1540), .S(n1514) );
  XNOR2_X1 U1595 ( .A(xmem_data[10]), .B(n1841), .ZN(n1498) );
  NOR2_X1 U1596 ( .A1(n1498), .A2(n1506), .ZN(n1505) );
  FA_X1 U1597 ( .A(n1505), .B(n1504), .CI(n1503), .CO(n1543), .S(n1539) );
  XNOR2_X1 U1598 ( .A(fmem_data[10]), .B(xmem_data[10]), .ZN(n1507) );
  OAI21_X1 U1599 ( .B1(n1221), .B2(n1219), .A(n1235), .ZN(n1508) );
  OR2_X1 U1600 ( .A1(n1543), .A2(n1542), .ZN(n1510) );
  NOR2_X1 U1601 ( .A1(n1509), .A2(n1219), .ZN(n1511) );
  AND2_X1 U1602 ( .A1(n1511), .A2(n1510), .ZN(n1914) );
  NAND2_X1 U1603 ( .A1(m_valid_y), .A2(m_ready_y), .ZN(n1945) );
  INV_X1 U1604 ( .A(reset), .ZN(n2407) );
  NAND2_X1 U1605 ( .A1(n1945), .A2(n2407), .ZN(n2379) );
  NOR2_X1 U1606 ( .A1(n2379), .A2(n2505), .ZN(n2381) );
  NOR2_X1 U1607 ( .A1(n2512), .A2(s_ready_x), .ZN(n1940) );
  NAND2_X1 U1608 ( .A1(n2381), .A2(n1940), .ZN(n1547) );
  BUF_X1 U1609 ( .A(n1216), .Z(n1601) );
  XNOR2_X1 U1610 ( .A(n1197), .B(n1528), .ZN(n1526) );
  NOR2_X1 U1611 ( .A1(n1526), .A2(n1224), .ZN(n1516) );
  INV_X1 U1612 ( .A(n1513), .ZN(n1515) );
  XNOR2_X1 U1613 ( .A(n1515), .B(n1514), .ZN(n1529) );
  INV_X1 U1614 ( .A(n1529), .ZN(n1532) );
  NOR2_X1 U1615 ( .A1(n1214), .A2(n1161), .ZN(n1535) );
  XOR2_X1 U1616 ( .A(n1518), .B(n1517), .Z(n1522) );
  NOR2_X1 U1617 ( .A1(n1522), .A2(n1521), .ZN(n1525) );
  NOR2_X1 U1618 ( .A1(n1525), .A2(n1519), .ZN(n1520) );
  NAND2_X1 U1619 ( .A1(n1535), .A2(n1520), .ZN(n1538) );
  NAND2_X1 U1620 ( .A1(n1522), .A2(n1521), .ZN(n1523) );
  OAI21_X1 U1621 ( .B1(n1525), .B2(n1524), .A(n1523), .ZN(n1536) );
  NAND2_X1 U1622 ( .A1(n1526), .A2(n1224), .ZN(n1533) );
  NAND2_X1 U1623 ( .A1(n1529), .A2(n1530), .ZN(n1531) );
  OAI21_X1 U1624 ( .B1(n1532), .B2(n1533), .A(n1531), .ZN(n1534) );
  AOI21_X1 U1625 ( .B1(n1536), .B2(n1215), .A(n1534), .ZN(n1537) );
  OAI21_X1 U1626 ( .B1(n1538), .B2(n1910), .A(n1537), .ZN(n1911) );
  HA_X1 U1627 ( .A(n1540), .B(n1539), .S(n1541) );
  INV_X1 U1628 ( .A(n1541), .ZN(n1546) );
  HA_X1 U1629 ( .A(n1543), .B(n1542), .S(n1544) );
  INV_X1 U1630 ( .A(n1544), .ZN(n1545) );
  NOR2_X1 U1631 ( .A1(n1546), .A2(n1545), .ZN(n1912) );
  OR2_X1 U1632 ( .A1(n1607), .A2(n1597), .ZN(n1553) );
  INV_X1 U1633 ( .A(n1549), .ZN(n1593) );
  OAI21_X1 U1634 ( .B1(n1550), .B2(n1593), .A(n1592), .ZN(n1606) );
  INV_X1 U1635 ( .A(n1606), .ZN(n1599) );
  OAI21_X1 U1636 ( .B1(n1607), .B2(n1603), .A(n1608), .ZN(n1551) );
  INV_X1 U1637 ( .A(n1551), .ZN(n1552) );
  OAI21_X1 U1638 ( .B1(n1553), .B2(n1599), .A(n1552), .ZN(n1554) );
  INV_X1 U1639 ( .A(n1940), .ZN(n1944) );
  NOR2_X1 U1640 ( .A1(n1920), .A2(n2507), .ZN(n1557) );
  AOI21_X1 U1641 ( .B1(n1213), .B2(n1558), .A(n1557), .ZN(n1559) );
  NAND2_X1 U1642 ( .A1(n1559), .A2(n1601), .ZN(n796) );
  AND2_X1 U1643 ( .A1(fmem_data[0]), .A2(xmem_data[0]), .ZN(n1560) );
  NAND2_X1 U1644 ( .A1(n1178), .A2(n1560), .ZN(n1563) );
  NAND3_X1 U1645 ( .A1(n1563), .A2(n1561), .A3(n1562), .ZN(n805) );
  OR2_X1 U1646 ( .A1(n1565), .A2(n1564), .ZN(n1567) );
  AND2_X1 U1647 ( .A1(n1567), .A2(n1566), .ZN(n1568) );
  NAND2_X1 U1648 ( .A1(n1178), .A2(n1568), .ZN(n1570) );
  NAND3_X1 U1649 ( .A1(n1570), .A2(n1561), .A3(n1569), .ZN(n804) );
  NAND2_X1 U1650 ( .A1(n1572), .A2(n1571), .ZN(n1574) );
  XNOR2_X1 U1651 ( .A(n1574), .B(n1573), .ZN(n1575) );
  NAND2_X1 U1652 ( .A1(n1178), .A2(n1575), .ZN(n1577) );
  NAND3_X1 U1653 ( .A1(n1577), .A2(n1561), .A3(n1576), .ZN(n803) );
  INV_X1 U1654 ( .A(n1578), .ZN(n1580) );
  NAND2_X1 U1655 ( .A1(n1580), .A2(n1579), .ZN(n1582) );
  XOR2_X1 U1656 ( .A(n1582), .B(n1581), .Z(n1583) );
  NAND2_X1 U1657 ( .A1(n1178), .A2(n1583), .ZN(n1585) );
  NAND3_X1 U1658 ( .A1(n1585), .A2(n1561), .A3(n1584), .ZN(n802) );
  INV_X1 U1659 ( .A(n1586), .ZN(n1588) );
  NAND2_X1 U1660 ( .A1(n1588), .A2(n1587), .ZN(n1589) );
  XOR2_X1 U1661 ( .A(n1589), .B(n1208), .Z(n1590) );
  NAND2_X1 U1662 ( .A1(n1213), .A2(n1590), .ZN(n1591) );
  NAND3_X1 U1663 ( .A1(n1591), .A2(n1601), .A3(n1240), .ZN(n800) );
  NAND2_X1 U1664 ( .A1(n1175), .A2(n1592), .ZN(n1594) );
  XOR2_X1 U1665 ( .A(n1594), .B(n1593), .Z(n1595) );
  NAND2_X1 U1666 ( .A1(n1178), .A2(n1595), .ZN(n1596) );
  NAND3_X1 U1667 ( .A1(n1596), .A2(n1601), .A3(n1241), .ZN(n799) );
  INV_X1 U1668 ( .A(n1597), .ZN(n1605) );
  NAND2_X1 U1669 ( .A1(n1605), .A2(n1603), .ZN(n1598) );
  XOR2_X1 U1670 ( .A(n1599), .B(n1598), .Z(n1600) );
  NAND2_X1 U1671 ( .A1(n1213), .A2(n1600), .ZN(n1602) );
  NAND3_X1 U1672 ( .A1(n1602), .A2(n1601), .A3(n1242), .ZN(n798) );
  INV_X1 U1673 ( .A(n1603), .ZN(n1604) );
  AOI21_X1 U1674 ( .B1(n1606), .B2(n1605), .A(n1604), .ZN(n1611) );
  INV_X1 U1675 ( .A(n1607), .ZN(n1609) );
  NAND2_X1 U1676 ( .A1(n1609), .A2(n1608), .ZN(n1610) );
  XOR2_X1 U1677 ( .A(n1611), .B(n1610), .Z(n1612) );
  NAND2_X1 U1678 ( .A1(n1213), .A2(n1612), .ZN(n1613) );
  NAND3_X1 U1679 ( .A1(n1613), .A2(n1561), .A3(n1243), .ZN(n797) );
  NAND2_X1 U1680 ( .A1(xmem_addr[3]), .A2(xmem_addr[4]), .ZN(n1938) );
  NAND2_X1 U1681 ( .A1(n2502), .A2(xmem_addr[2]), .ZN(n1952) );
  INV_X1 U1682 ( .A(n1952), .ZN(n1614) );
  NAND2_X1 U1683 ( .A1(n1614), .A2(n2493), .ZN(n2346) );
  NOR2_X1 U1684 ( .A1(n1938), .A2(n2346), .ZN(n1871) );
  NAND2_X1 U1685 ( .A1(xmem_addr[0]), .A2(n1614), .ZN(n2247) );
  NOR2_X1 U1686 ( .A1(n2247), .A2(n1938), .ZN(n1870) );
  AOI22_X1 U1687 ( .A1(n1871), .A2(\xmem_inst/mem[28][6] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][6] ), .ZN(n1618) );
  NOR2_X1 U1688 ( .A1(xmem_addr[3]), .A2(xmem_addr[4]), .ZN(n1963) );
  NAND2_X1 U1689 ( .A1(n1963), .A2(n2493), .ZN(n1626) );
  NOR2_X1 U1690 ( .A1(n1952), .A2(n1626), .ZN(n1873) );
  NOR2_X1 U1691 ( .A1(xmem_addr[4]), .A2(n2495), .ZN(n2071) );
  NAND2_X1 U1692 ( .A1(n2071), .A2(n2493), .ZN(n1627) );
  NOR2_X1 U1693 ( .A1(n1952), .A2(n1627), .ZN(n1872) );
  AOI22_X1 U1694 ( .A1(n1873), .A2(\xmem_inst/mem[4][6] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][6] ), .ZN(n1617) );
  NAND2_X1 U1695 ( .A1(xmem_addr[1]), .A2(xmem_addr[2]), .ZN(n1634) );
  NOR2_X1 U1696 ( .A1(n1634), .A2(n1627), .ZN(n2151) );
  NOR2_X1 U1697 ( .A1(n1634), .A2(n1626), .ZN(n2043) );
  AOI22_X1 U1698 ( .A1(n2151), .A2(\xmem_inst/mem[14][6] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][6] ), .ZN(n1616) );
  NAND2_X1 U1699 ( .A1(xmem_addr[4]), .A2(n2495), .ZN(n1961) );
  NOR2_X1 U1700 ( .A1(n1961), .A2(n2346), .ZN(n1875) );
  NOR2_X1 U1701 ( .A1(n2247), .A2(n1961), .ZN(n1874) );
  AOI22_X1 U1702 ( .A1(n1875), .A2(\xmem_inst/mem[20][6] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][6] ), .ZN(n1615) );
  NAND4_X1 U1703 ( .A1(n1618), .A2(n1617), .A3(n1616), .A4(n1615), .ZN(n1643)
         );
  NOR2_X1 U1704 ( .A1(xmem_addr[2]), .A2(n2502), .ZN(n1619) );
  NAND2_X1 U1705 ( .A1(n1619), .A2(n2493), .ZN(n2318) );
  NOR2_X1 U1706 ( .A1(n1938), .A2(n2318), .ZN(n1859) );
  INV_X1 U1707 ( .A(n1619), .ZN(n1620) );
  NOR2_X1 U1708 ( .A1(n1620), .A2(n1627), .ZN(n1858) );
  AOI22_X1 U1709 ( .A1(n1859), .A2(\xmem_inst/mem[26][6] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][6] ), .ZN(n1624) );
  NOR2_X1 U1710 ( .A1(n1620), .A2(n1626), .ZN(n1861) );
  NAND2_X1 U1711 ( .A1(xmem_addr[0]), .A2(n1619), .ZN(n2332) );
  NOR2_X1 U1712 ( .A1(n1938), .A2(n2332), .ZN(n1860) );
  AOI22_X1 U1713 ( .A1(n1861), .A2(\xmem_inst/mem[2][6] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][6] ), .ZN(n1623) );
  NOR2_X1 U1714 ( .A1(n1961), .A2(n2318), .ZN(n1863) );
  NAND2_X1 U1715 ( .A1(xmem_addr[0]), .A2(n1963), .ZN(n1633) );
  NOR2_X1 U1716 ( .A1(n1620), .A2(n1633), .ZN(n1862) );
  AOI22_X1 U1717 ( .A1(n1863), .A2(\xmem_inst/mem[18][6] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][6] ), .ZN(n1622) );
  NAND2_X1 U1718 ( .A1(xmem_addr[0]), .A2(n2071), .ZN(n1635) );
  NOR2_X1 U1719 ( .A1(n1620), .A2(n1635), .ZN(n1865) );
  NOR2_X1 U1720 ( .A1(n2332), .A2(n1961), .ZN(n1864) );
  AOI22_X1 U1721 ( .A1(n1865), .A2(\xmem_inst/mem[11][6] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][6] ), .ZN(n1621) );
  NAND4_X1 U1722 ( .A1(n1624), .A2(n1623), .A3(n1622), .A4(n1621), .ZN(n1642)
         );
  NOR2_X1 U1723 ( .A1(xmem_addr[1]), .A2(xmem_addr[2]), .ZN(n1625) );
  NAND2_X1 U1724 ( .A1(n1625), .A2(n2493), .ZN(n2290) );
  NOR2_X1 U1725 ( .A1(n1938), .A2(n2290), .ZN(n1847) );
  NAND2_X1 U1726 ( .A1(xmem_addr[0]), .A2(n1625), .ZN(n2304) );
  NOR2_X1 U1727 ( .A1(n1938), .A2(n2304), .ZN(n1846) );
  AOI22_X1 U1728 ( .A1(n1847), .A2(\xmem_inst/mem[24][6] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][6] ), .ZN(n1632) );
  INV_X1 U1729 ( .A(n1625), .ZN(n1628) );
  NOR2_X1 U1730 ( .A1(n1628), .A2(n1626), .ZN(n1849) );
  NOR2_X1 U1731 ( .A1(n1628), .A2(n1627), .ZN(n1848) );
  AOI22_X1 U1732 ( .A1(n1849), .A2(\xmem_inst/mem[0][6] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][6] ), .ZN(n1631) );
  NOR2_X1 U1733 ( .A1(n1961), .A2(n2290), .ZN(n1851) );
  NOR2_X1 U1734 ( .A1(n1633), .A2(n1628), .ZN(n1850) );
  AOI22_X1 U1735 ( .A1(n1851), .A2(\xmem_inst/mem[16][6] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][6] ), .ZN(n1630) );
  NOR2_X1 U1736 ( .A1(n1635), .A2(n1628), .ZN(n1853) );
  NOR2_X1 U1737 ( .A1(n1961), .A2(n2304), .ZN(n1852) );
  AOI22_X1 U1738 ( .A1(n1853), .A2(\xmem_inst/mem[9][6] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][6] ), .ZN(n1629) );
  NAND4_X1 U1739 ( .A1(n1632), .A2(n1631), .A3(n1630), .A4(n1629), .ZN(n1641)
         );
  NOR3_X2 U1740 ( .A1(xmem_addr[0]), .A2(n1634), .A3(n1961), .ZN(n2261) );
  NAND2_X1 U1741 ( .A1(n2261), .A2(\xmem_inst/mem[22][6] ), .ZN(n1639) );
  NOR2_X1 U1742 ( .A1(n1634), .A2(n1633), .ZN(n2057) );
  NOR2_X1 U1743 ( .A1(n1952), .A2(n1633), .ZN(n1884) );
  AOI22_X1 U1744 ( .A1(n2057), .A2(\xmem_inst/mem[7][6] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][6] ), .ZN(n1638) );
  NOR2_X1 U1745 ( .A1(n2493), .A2(n1634), .ZN(n1955) );
  NAND2_X1 U1746 ( .A1(n1955), .A2(n2071), .ZN(n2165) );
  INV_X1 U1747 ( .A(n2165), .ZN(n1885) );
  INV_X1 U1748 ( .A(n1961), .ZN(n2180) );
  AND2_X1 U1749 ( .A1(n1955), .A2(n2180), .ZN(n2275) );
  AOI22_X1 U1750 ( .A1(\xmem_inst/mem[15][6] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][6] ), .ZN(n1637) );
  NOR2_X1 U1751 ( .A1(n1952), .A2(n1635), .ZN(n1883) );
  NAND2_X1 U1752 ( .A1(n1883), .A2(\xmem_inst/mem[13][6] ), .ZN(n1636) );
  NAND4_X1 U1753 ( .A1(n1639), .A2(n1638), .A3(n1637), .A4(n1636), .ZN(n1640)
         );
  AOI22_X1 U1754 ( .A1(n1871), .A2(\xmem_inst/mem[28][0] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][0] ), .ZN(n1647) );
  AOI22_X1 U1755 ( .A1(n1873), .A2(\xmem_inst/mem[4][0] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][0] ), .ZN(n1646) );
  AOI22_X1 U1756 ( .A1(n2151), .A2(\xmem_inst/mem[14][0] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][0] ), .ZN(n1645) );
  AOI22_X1 U1757 ( .A1(n1875), .A2(\xmem_inst/mem[20][0] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][0] ), .ZN(n1644) );
  NAND4_X1 U1758 ( .A1(n1647), .A2(n1646), .A3(n1645), .A4(n1644), .ZN(n1663)
         );
  AOI22_X1 U1759 ( .A1(n1859), .A2(\xmem_inst/mem[26][0] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][0] ), .ZN(n1651) );
  AOI22_X1 U1760 ( .A1(n1861), .A2(\xmem_inst/mem[2][0] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][0] ), .ZN(n1650) );
  AOI22_X1 U1761 ( .A1(n1863), .A2(\xmem_inst/mem[18][0] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][0] ), .ZN(n1649) );
  AOI22_X1 U1762 ( .A1(n1865), .A2(\xmem_inst/mem[11][0] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][0] ), .ZN(n1648) );
  NAND4_X1 U1763 ( .A1(n1651), .A2(n1650), .A3(n1649), .A4(n1648), .ZN(n1662)
         );
  AOI22_X1 U1764 ( .A1(n1847), .A2(\xmem_inst/mem[24][0] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][0] ), .ZN(n1655) );
  AOI22_X1 U1765 ( .A1(n1849), .A2(\xmem_inst/mem[0][0] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][0] ), .ZN(n1654) );
  AOI22_X1 U1766 ( .A1(n1851), .A2(\xmem_inst/mem[16][0] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][0] ), .ZN(n1653) );
  AOI22_X1 U1767 ( .A1(n1853), .A2(\xmem_inst/mem[9][0] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][0] ), .ZN(n1652) );
  NAND4_X1 U1768 ( .A1(n1655), .A2(n1654), .A3(n1653), .A4(n1652), .ZN(n1661)
         );
  NAND2_X1 U1769 ( .A1(n2261), .A2(\xmem_inst/mem[22][0] ), .ZN(n1659) );
  AOI22_X1 U1770 ( .A1(n2057), .A2(\xmem_inst/mem[7][0] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][0] ), .ZN(n1658) );
  AOI22_X1 U1771 ( .A1(\xmem_inst/mem[15][0] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][0] ), .ZN(n1657) );
  NAND2_X1 U1772 ( .A1(n1883), .A2(\xmem_inst/mem[13][0] ), .ZN(n1656) );
  NAND4_X1 U1773 ( .A1(n1659), .A2(n1658), .A3(n1657), .A4(n1656), .ZN(n1660)
         );
  AOI22_X1 U1774 ( .A1(n1871), .A2(\xmem_inst/mem[28][1] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][1] ), .ZN(n1667) );
  AOI22_X1 U1775 ( .A1(n1873), .A2(\xmem_inst/mem[4][1] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][1] ), .ZN(n1666) );
  AOI22_X1 U1776 ( .A1(n2151), .A2(\xmem_inst/mem[14][1] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][1] ), .ZN(n1665) );
  AOI22_X1 U1777 ( .A1(n1875), .A2(\xmem_inst/mem[20][1] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][1] ), .ZN(n1664) );
  NAND4_X1 U1778 ( .A1(n1667), .A2(n1666), .A3(n1665), .A4(n1664), .ZN(n1683)
         );
  AOI22_X1 U1779 ( .A1(n1859), .A2(\xmem_inst/mem[26][1] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][1] ), .ZN(n1671) );
  AOI22_X1 U1780 ( .A1(n1861), .A2(\xmem_inst/mem[2][1] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][1] ), .ZN(n1670) );
  AOI22_X1 U1781 ( .A1(n1863), .A2(\xmem_inst/mem[18][1] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][1] ), .ZN(n1669) );
  AOI22_X1 U1782 ( .A1(n1865), .A2(\xmem_inst/mem[11][1] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][1] ), .ZN(n1668) );
  NAND4_X1 U1783 ( .A1(n1671), .A2(n1670), .A3(n1669), .A4(n1668), .ZN(n1682)
         );
  AOI22_X1 U1784 ( .A1(n1847), .A2(\xmem_inst/mem[24][1] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][1] ), .ZN(n1675) );
  AOI22_X1 U1785 ( .A1(n1849), .A2(\xmem_inst/mem[0][1] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][1] ), .ZN(n1674) );
  AOI22_X1 U1786 ( .A1(n1851), .A2(\xmem_inst/mem[16][1] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][1] ), .ZN(n1673) );
  AOI22_X1 U1787 ( .A1(n1853), .A2(\xmem_inst/mem[9][1] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][1] ), .ZN(n1672) );
  NAND4_X1 U1788 ( .A1(n1675), .A2(n1674), .A3(n1673), .A4(n1672), .ZN(n1681)
         );
  NAND2_X1 U1789 ( .A1(n2261), .A2(\xmem_inst/mem[22][1] ), .ZN(n1679) );
  AOI22_X1 U1790 ( .A1(n2057), .A2(\xmem_inst/mem[7][1] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][1] ), .ZN(n1678) );
  AOI22_X1 U1791 ( .A1(\xmem_inst/mem[15][1] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][1] ), .ZN(n1677) );
  NAND2_X1 U1792 ( .A1(n1883), .A2(\xmem_inst/mem[13][1] ), .ZN(n1676) );
  NAND4_X1 U1793 ( .A1(n1679), .A2(n1678), .A3(n1677), .A4(n1676), .ZN(n1680)
         );
  AOI22_X1 U1794 ( .A1(n1871), .A2(\xmem_inst/mem[28][9] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][9] ), .ZN(n1687) );
  AOI22_X1 U1795 ( .A1(n1873), .A2(\xmem_inst/mem[4][9] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][9] ), .ZN(n1686) );
  AOI22_X1 U1796 ( .A1(n2151), .A2(\xmem_inst/mem[14][9] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][9] ), .ZN(n1685) );
  AOI22_X1 U1797 ( .A1(n1875), .A2(\xmem_inst/mem[20][9] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][9] ), .ZN(n1684) );
  NAND4_X1 U1798 ( .A1(n1687), .A2(n1686), .A3(n1685), .A4(n1684), .ZN(n1703)
         );
  AOI22_X1 U1799 ( .A1(n1859), .A2(\xmem_inst/mem[26][9] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][9] ), .ZN(n1691) );
  AOI22_X1 U1800 ( .A1(n1861), .A2(\xmem_inst/mem[2][9] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][9] ), .ZN(n1690) );
  AOI22_X1 U1801 ( .A1(n1863), .A2(\xmem_inst/mem[18][9] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][9] ), .ZN(n1689) );
  AOI22_X1 U1802 ( .A1(n1865), .A2(\xmem_inst/mem[11][9] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][9] ), .ZN(n1688) );
  NAND4_X1 U1803 ( .A1(n1691), .A2(n1690), .A3(n1689), .A4(n1688), .ZN(n1702)
         );
  AOI22_X1 U1804 ( .A1(n1847), .A2(\xmem_inst/mem[24][9] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][9] ), .ZN(n1695) );
  AOI22_X1 U1805 ( .A1(n1849), .A2(\xmem_inst/mem[0][9] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][9] ), .ZN(n1694) );
  AOI22_X1 U1806 ( .A1(n1851), .A2(\xmem_inst/mem[16][9] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][9] ), .ZN(n1693) );
  AOI22_X1 U1807 ( .A1(n1853), .A2(\xmem_inst/mem[9][9] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][9] ), .ZN(n1692) );
  NAND4_X1 U1808 ( .A1(n1695), .A2(n1694), .A3(n1693), .A4(n1692), .ZN(n1701)
         );
  NAND2_X1 U1809 ( .A1(n2261), .A2(\xmem_inst/mem[22][9] ), .ZN(n1699) );
  AOI22_X1 U1810 ( .A1(n2057), .A2(\xmem_inst/mem[7][9] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][9] ), .ZN(n1698) );
  AOI22_X1 U1811 ( .A1(\xmem_inst/mem[15][9] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][9] ), .ZN(n1697) );
  NAND2_X1 U1812 ( .A1(n1883), .A2(\xmem_inst/mem[13][9] ), .ZN(n1696) );
  NAND4_X1 U1813 ( .A1(n1699), .A2(n1698), .A3(n1697), .A4(n1696), .ZN(n1700)
         );
  AOI22_X1 U1814 ( .A1(n1871), .A2(\xmem_inst/mem[28][5] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][5] ), .ZN(n1707) );
  AOI22_X1 U1815 ( .A1(n1873), .A2(\xmem_inst/mem[4][5] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][5] ), .ZN(n1706) );
  AOI22_X1 U1816 ( .A1(n2151), .A2(\xmem_inst/mem[14][5] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][5] ), .ZN(n1705) );
  AOI22_X1 U1817 ( .A1(n1875), .A2(\xmem_inst/mem[20][5] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][5] ), .ZN(n1704) );
  NAND4_X1 U1818 ( .A1(n1707), .A2(n1706), .A3(n1705), .A4(n1704), .ZN(n1723)
         );
  AOI22_X1 U1819 ( .A1(n1859), .A2(\xmem_inst/mem[26][5] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][5] ), .ZN(n1711) );
  AOI22_X1 U1820 ( .A1(n1861), .A2(\xmem_inst/mem[2][5] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][5] ), .ZN(n1710) );
  AOI22_X1 U1821 ( .A1(n1863), .A2(\xmem_inst/mem[18][5] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][5] ), .ZN(n1709) );
  AOI22_X1 U1822 ( .A1(n1865), .A2(\xmem_inst/mem[11][5] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][5] ), .ZN(n1708) );
  NAND4_X1 U1823 ( .A1(n1711), .A2(n1710), .A3(n1709), .A4(n1708), .ZN(n1722)
         );
  AOI22_X1 U1824 ( .A1(n1847), .A2(\xmem_inst/mem[24][5] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][5] ), .ZN(n1715) );
  AOI22_X1 U1825 ( .A1(n1849), .A2(\xmem_inst/mem[0][5] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][5] ), .ZN(n1714) );
  AOI22_X1 U1826 ( .A1(n1851), .A2(\xmem_inst/mem[16][5] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][5] ), .ZN(n1713) );
  AOI22_X1 U1827 ( .A1(n1853), .A2(\xmem_inst/mem[9][5] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][5] ), .ZN(n1712) );
  NAND4_X1 U1828 ( .A1(n1715), .A2(n1714), .A3(n1713), .A4(n1712), .ZN(n1721)
         );
  NAND2_X1 U1829 ( .A1(n2261), .A2(\xmem_inst/mem[22][5] ), .ZN(n1719) );
  AOI22_X1 U1830 ( .A1(n2057), .A2(\xmem_inst/mem[7][5] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][5] ), .ZN(n1718) );
  AOI22_X1 U1831 ( .A1(\xmem_inst/mem[15][5] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][5] ), .ZN(n1717) );
  NAND2_X1 U1832 ( .A1(n1883), .A2(\xmem_inst/mem[13][5] ), .ZN(n1716) );
  NAND4_X1 U1833 ( .A1(n1719), .A2(n1718), .A3(n1717), .A4(n1716), .ZN(n1720)
         );
  AOI22_X1 U1834 ( .A1(n1871), .A2(\xmem_inst/mem[28][3] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][3] ), .ZN(n1727) );
  AOI22_X1 U1835 ( .A1(n1873), .A2(\xmem_inst/mem[4][3] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][3] ), .ZN(n1726) );
  AOI22_X1 U1836 ( .A1(n2151), .A2(\xmem_inst/mem[14][3] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][3] ), .ZN(n1725) );
  AOI22_X1 U1837 ( .A1(n1875), .A2(\xmem_inst/mem[20][3] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][3] ), .ZN(n1724) );
  NAND4_X1 U1838 ( .A1(n1727), .A2(n1726), .A3(n1725), .A4(n1724), .ZN(n1743)
         );
  AOI22_X1 U1839 ( .A1(n1859), .A2(\xmem_inst/mem[26][3] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][3] ), .ZN(n1731) );
  AOI22_X1 U1840 ( .A1(n1861), .A2(\xmem_inst/mem[2][3] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][3] ), .ZN(n1730) );
  AOI22_X1 U1841 ( .A1(n1863), .A2(\xmem_inst/mem[18][3] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][3] ), .ZN(n1729) );
  AOI22_X1 U1842 ( .A1(n1865), .A2(\xmem_inst/mem[11][3] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][3] ), .ZN(n1728) );
  NAND4_X1 U1843 ( .A1(n1731), .A2(n1730), .A3(n1729), .A4(n1728), .ZN(n1742)
         );
  AOI22_X1 U1844 ( .A1(n1847), .A2(\xmem_inst/mem[24][3] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][3] ), .ZN(n1735) );
  AOI22_X1 U1845 ( .A1(n1849), .A2(\xmem_inst/mem[0][3] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][3] ), .ZN(n1734) );
  AOI22_X1 U1846 ( .A1(n1851), .A2(\xmem_inst/mem[16][3] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][3] ), .ZN(n1733) );
  AOI22_X1 U1847 ( .A1(n1853), .A2(\xmem_inst/mem[9][3] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][3] ), .ZN(n1732) );
  NAND4_X1 U1848 ( .A1(n1735), .A2(n1734), .A3(n1733), .A4(n1732), .ZN(n1741)
         );
  NAND2_X1 U1849 ( .A1(n2261), .A2(\xmem_inst/mem[22][3] ), .ZN(n1739) );
  AOI22_X1 U1850 ( .A1(n2057), .A2(\xmem_inst/mem[7][3] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][3] ), .ZN(n1738) );
  AOI22_X1 U1851 ( .A1(\xmem_inst/mem[15][3] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][3] ), .ZN(n1737) );
  NAND2_X1 U1852 ( .A1(n1883), .A2(\xmem_inst/mem[13][3] ), .ZN(n1736) );
  NAND4_X1 U1853 ( .A1(n1739), .A2(n1738), .A3(n1737), .A4(n1736), .ZN(n1740)
         );
  NAND2_X1 U1854 ( .A1(n1745), .A2(n1744), .ZN(n1747) );
  XNOR2_X1 U1855 ( .A(n1747), .B(n1746), .ZN(n1748) );
  NAND2_X1 U1856 ( .A1(n1178), .A2(n1748), .ZN(n1753) );
  OAI21_X1 U1857 ( .B1(n1164), .B2(n1248), .A(n1751), .ZN(n1752) );
  NAND2_X1 U1858 ( .A1(n1753), .A2(n1752), .ZN(n801) );
  AOI22_X1 U1859 ( .A1(n1871), .A2(\xmem_inst/mem[28][4] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][4] ), .ZN(n1757) );
  AOI22_X1 U1860 ( .A1(n1873), .A2(\xmem_inst/mem[4][4] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][4] ), .ZN(n1756) );
  AOI22_X1 U1861 ( .A1(n2151), .A2(\xmem_inst/mem[14][4] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][4] ), .ZN(n1755) );
  AOI22_X1 U1862 ( .A1(n1875), .A2(\xmem_inst/mem[20][4] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][4] ), .ZN(n1754) );
  NAND4_X1 U1863 ( .A1(n1757), .A2(n1756), .A3(n1755), .A4(n1754), .ZN(n1773)
         );
  AOI22_X1 U1864 ( .A1(n1859), .A2(\xmem_inst/mem[26][4] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][4] ), .ZN(n1761) );
  AOI22_X1 U1865 ( .A1(n1861), .A2(\xmem_inst/mem[2][4] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][4] ), .ZN(n1760) );
  AOI22_X1 U1866 ( .A1(n1863), .A2(\xmem_inst/mem[18][4] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][4] ), .ZN(n1759) );
  AOI22_X1 U1867 ( .A1(n1865), .A2(\xmem_inst/mem[11][4] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][4] ), .ZN(n1758) );
  NAND4_X1 U1868 ( .A1(n1761), .A2(n1760), .A3(n1759), .A4(n1758), .ZN(n1772)
         );
  AOI22_X1 U1869 ( .A1(n1847), .A2(\xmem_inst/mem[24][4] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][4] ), .ZN(n1765) );
  AOI22_X1 U1870 ( .A1(n1849), .A2(\xmem_inst/mem[0][4] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][4] ), .ZN(n1764) );
  AOI22_X1 U1871 ( .A1(n1851), .A2(\xmem_inst/mem[16][4] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][4] ), .ZN(n1763) );
  AOI22_X1 U1872 ( .A1(n1853), .A2(\xmem_inst/mem[9][4] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][4] ), .ZN(n1762) );
  NAND4_X1 U1873 ( .A1(n1765), .A2(n1764), .A3(n1763), .A4(n1762), .ZN(n1771)
         );
  NAND2_X1 U1874 ( .A1(n2261), .A2(\xmem_inst/mem[22][4] ), .ZN(n1769) );
  AOI22_X1 U1875 ( .A1(n2057), .A2(\xmem_inst/mem[7][4] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][4] ), .ZN(n1768) );
  AOI22_X1 U1876 ( .A1(\xmem_inst/mem[15][4] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][4] ), .ZN(n1767) );
  NAND2_X1 U1877 ( .A1(n1883), .A2(\xmem_inst/mem[13][4] ), .ZN(n1766) );
  NAND4_X1 U1878 ( .A1(n1769), .A2(n1768), .A3(n1767), .A4(n1766), .ZN(n1770)
         );
  OR4_X1 U1879 ( .A1(n1773), .A2(n1772), .A3(n1771), .A4(n1770), .ZN(
        \xmem_inst/N22 ) );
  AOI22_X1 U1880 ( .A1(n1871), .A2(\xmem_inst/mem[28][2] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][2] ), .ZN(n1777) );
  AOI22_X1 U1881 ( .A1(n1873), .A2(\xmem_inst/mem[4][2] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][2] ), .ZN(n1776) );
  AOI22_X1 U1882 ( .A1(n2151), .A2(\xmem_inst/mem[14][2] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][2] ), .ZN(n1775) );
  AOI22_X1 U1883 ( .A1(n1875), .A2(\xmem_inst/mem[20][2] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][2] ), .ZN(n1774) );
  NAND4_X1 U1884 ( .A1(n1777), .A2(n1776), .A3(n1775), .A4(n1774), .ZN(n1793)
         );
  AOI22_X1 U1885 ( .A1(n1859), .A2(\xmem_inst/mem[26][2] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][2] ), .ZN(n1781) );
  AOI22_X1 U1886 ( .A1(n1861), .A2(\xmem_inst/mem[2][2] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][2] ), .ZN(n1780) );
  AOI22_X1 U1887 ( .A1(n1863), .A2(\xmem_inst/mem[18][2] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][2] ), .ZN(n1779) );
  AOI22_X1 U1888 ( .A1(n1865), .A2(\xmem_inst/mem[11][2] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][2] ), .ZN(n1778) );
  NAND4_X1 U1889 ( .A1(n1781), .A2(n1780), .A3(n1779), .A4(n1778), .ZN(n1792)
         );
  AOI22_X1 U1890 ( .A1(n1847), .A2(\xmem_inst/mem[24][2] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][2] ), .ZN(n1785) );
  AOI22_X1 U1891 ( .A1(n1849), .A2(\xmem_inst/mem[0][2] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][2] ), .ZN(n1784) );
  AOI22_X1 U1892 ( .A1(n1851), .A2(\xmem_inst/mem[16][2] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][2] ), .ZN(n1783) );
  AOI22_X1 U1893 ( .A1(n1853), .A2(\xmem_inst/mem[9][2] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][2] ), .ZN(n1782) );
  NAND4_X1 U1894 ( .A1(n1785), .A2(n1784), .A3(n1783), .A4(n1782), .ZN(n1791)
         );
  NAND2_X1 U1895 ( .A1(n2261), .A2(\xmem_inst/mem[22][2] ), .ZN(n1789) );
  AOI22_X1 U1896 ( .A1(n2057), .A2(\xmem_inst/mem[7][2] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][2] ), .ZN(n1788) );
  AOI22_X1 U1897 ( .A1(\xmem_inst/mem[15][2] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][2] ), .ZN(n1787) );
  NAND2_X1 U1898 ( .A1(n1883), .A2(\xmem_inst/mem[13][2] ), .ZN(n1786) );
  NAND4_X1 U1899 ( .A1(n1789), .A2(n1788), .A3(n1787), .A4(n1786), .ZN(n1790)
         );
  OR4_X1 U1900 ( .A1(n1793), .A2(n1792), .A3(n1791), .A4(n1790), .ZN(
        \xmem_inst/N24 ) );
  AOI22_X1 U1901 ( .A1(n1871), .A2(\xmem_inst/mem[28][8] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][8] ), .ZN(n1797) );
  AOI22_X1 U1902 ( .A1(n1873), .A2(\xmem_inst/mem[4][8] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][8] ), .ZN(n1796) );
  AOI22_X1 U1903 ( .A1(n2151), .A2(\xmem_inst/mem[14][8] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][8] ), .ZN(n1795) );
  AOI22_X1 U1904 ( .A1(n1875), .A2(\xmem_inst/mem[20][8] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][8] ), .ZN(n1794) );
  NAND4_X1 U1905 ( .A1(n1797), .A2(n1796), .A3(n1795), .A4(n1794), .ZN(n1813)
         );
  AOI22_X1 U1906 ( .A1(n1859), .A2(\xmem_inst/mem[26][8] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][8] ), .ZN(n1801) );
  AOI22_X1 U1907 ( .A1(n1861), .A2(\xmem_inst/mem[2][8] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][8] ), .ZN(n1800) );
  AOI22_X1 U1908 ( .A1(n1863), .A2(\xmem_inst/mem[18][8] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][8] ), .ZN(n1799) );
  AOI22_X1 U1909 ( .A1(n1865), .A2(\xmem_inst/mem[11][8] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][8] ), .ZN(n1798) );
  NAND4_X1 U1910 ( .A1(n1801), .A2(n1800), .A3(n1799), .A4(n1798), .ZN(n1812)
         );
  AOI22_X1 U1911 ( .A1(n1847), .A2(\xmem_inst/mem[24][8] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][8] ), .ZN(n1805) );
  AOI22_X1 U1912 ( .A1(n1849), .A2(\xmem_inst/mem[0][8] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][8] ), .ZN(n1804) );
  AOI22_X1 U1913 ( .A1(n1851), .A2(\xmem_inst/mem[16][8] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][8] ), .ZN(n1803) );
  AOI22_X1 U1914 ( .A1(n1853), .A2(\xmem_inst/mem[9][8] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][8] ), .ZN(n1802) );
  NAND4_X1 U1915 ( .A1(n1805), .A2(n1804), .A3(n1803), .A4(n1802), .ZN(n1811)
         );
  NAND2_X1 U1916 ( .A1(n2261), .A2(\xmem_inst/mem[22][8] ), .ZN(n1809) );
  AOI22_X1 U1917 ( .A1(n2057), .A2(\xmem_inst/mem[7][8] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][8] ), .ZN(n1808) );
  AOI22_X1 U1918 ( .A1(\xmem_inst/mem[15][8] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][8] ), .ZN(n1807) );
  NAND2_X1 U1919 ( .A1(n1883), .A2(\xmem_inst/mem[13][8] ), .ZN(n1806) );
  NAND4_X1 U1920 ( .A1(n1809), .A2(n1808), .A3(n1807), .A4(n1806), .ZN(n1810)
         );
  OR4_X1 U1921 ( .A1(n1813), .A2(n1812), .A3(n1811), .A4(n1810), .ZN(
        \xmem_inst/N18 ) );
  AOI22_X1 U1922 ( .A1(n1871), .A2(\xmem_inst/mem[28][7] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][7] ), .ZN(n1817) );
  AOI22_X1 U1923 ( .A1(n1873), .A2(\xmem_inst/mem[4][7] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][7] ), .ZN(n1816) );
  AOI22_X1 U1924 ( .A1(n2151), .A2(\xmem_inst/mem[14][7] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][7] ), .ZN(n1815) );
  AOI22_X1 U1925 ( .A1(n1875), .A2(\xmem_inst/mem[20][7] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][7] ), .ZN(n1814) );
  NAND4_X1 U1926 ( .A1(n1817), .A2(n1816), .A3(n1815), .A4(n1814), .ZN(n1833)
         );
  AOI22_X1 U1927 ( .A1(n1859), .A2(\xmem_inst/mem[26][7] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][7] ), .ZN(n1821) );
  AOI22_X1 U1928 ( .A1(n1861), .A2(\xmem_inst/mem[2][7] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][7] ), .ZN(n1820) );
  AOI22_X1 U1929 ( .A1(n1863), .A2(\xmem_inst/mem[18][7] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][7] ), .ZN(n1819) );
  AOI22_X1 U1930 ( .A1(n1865), .A2(\xmem_inst/mem[11][7] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][7] ), .ZN(n1818) );
  NAND4_X1 U1931 ( .A1(n1821), .A2(n1820), .A3(n1819), .A4(n1818), .ZN(n1832)
         );
  AOI22_X1 U1932 ( .A1(n1847), .A2(\xmem_inst/mem[24][7] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][7] ), .ZN(n1825) );
  AOI22_X1 U1933 ( .A1(n1849), .A2(\xmem_inst/mem[0][7] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][7] ), .ZN(n1824) );
  AOI22_X1 U1934 ( .A1(n1851), .A2(\xmem_inst/mem[16][7] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][7] ), .ZN(n1823) );
  AOI22_X1 U1935 ( .A1(n1853), .A2(\xmem_inst/mem[9][7] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][7] ), .ZN(n1822) );
  NAND4_X1 U1936 ( .A1(n1825), .A2(n1824), .A3(n1823), .A4(n1822), .ZN(n1831)
         );
  NAND2_X1 U1937 ( .A1(n2261), .A2(\xmem_inst/mem[22][7] ), .ZN(n1829) );
  AOI22_X1 U1938 ( .A1(n2057), .A2(\xmem_inst/mem[7][7] ), .B1(n1884), .B2(
        \xmem_inst/mem[5][7] ), .ZN(n1828) );
  AOI22_X1 U1939 ( .A1(\xmem_inst/mem[15][7] ), .A2(n1885), .B1(n2275), .B2(
        \xmem_inst/mem[23][7] ), .ZN(n1827) );
  NAND2_X1 U1940 ( .A1(n1883), .A2(\xmem_inst/mem[13][7] ), .ZN(n1826) );
  NAND4_X1 U1941 ( .A1(n1829), .A2(n1828), .A3(n1827), .A4(n1826), .ZN(n1830)
         );
  OR4_X1 U1942 ( .A1(n1833), .A2(n1832), .A3(n1831), .A4(n1830), .ZN(
        \xmem_inst/N19 ) );
  NOR2_X1 U1943 ( .A1(fmem_addr[1]), .A2(fmem_addr[2]), .ZN(n1890) );
  NAND2_X1 U1944 ( .A1(n1890), .A2(n2496), .ZN(n1923) );
  NAND2_X1 U1945 ( .A1(n1923), .A2(fmem_addr[3]), .ZN(n1839) );
  NAND2_X1 U1946 ( .A1(n2496), .A2(fmem_addr[2]), .ZN(n1835) );
  NAND3_X1 U1947 ( .A1(n1923), .A2(n2498), .A3(n1835), .ZN(n1834) );
  OAI21_X1 U1948 ( .B1(n1839), .B2(n2500), .A(n1834), .ZN(n809) );
  OAI22_X1 U1949 ( .A1(n1839), .A2(n2499), .B1(fmem_addr[3]), .B2(n2491), .ZN(
        n811) );
  NAND2_X1 U1950 ( .A1(n2491), .A2(fmem_addr[0]), .ZN(n1894) );
  AOI22_X1 U1951 ( .A1(n1894), .A2(n1835), .B1(fmem_addr[2]), .B2(n2491), .ZN(
        n1836) );
  OAI22_X1 U1952 ( .A1(n1839), .A2(n2494), .B1(n1836), .B2(fmem_addr[3]), .ZN(
        n812) );
  NOR3_X1 U1953 ( .A1(n2491), .A2(fmem_addr[0]), .A3(n2489), .ZN(n1838) );
  INV_X1 U1954 ( .A(n1894), .ZN(n1837) );
  AOI211_X1 U1955 ( .C1(fmem_addr[0]), .C2(n2489), .A(n1838), .B(n1837), .ZN(
        n1840) );
  OAI22_X1 U1956 ( .A1(n1840), .A2(fmem_addr[3]), .B1(n1839), .B2(n2504), .ZN(
        n807) );
  INV_X1 U1957 ( .A(n1890), .ZN(n1843) );
  INV_X1 U1958 ( .A(n1923), .ZN(n1845) );
  OAI21_X1 U1959 ( .B1(n1845), .B2(n1841), .A(fmem_addr[3]), .ZN(n1842) );
  OAI21_X1 U1960 ( .B1(fmem_addr[3]), .B2(n1843), .A(n1842), .ZN(n808) );
  NAND2_X1 U1961 ( .A1(fmem_addr[0]), .A2(fmem_addr[2]), .ZN(n1844) );
  NOR2_X1 U1962 ( .A1(n1844), .A2(fmem_addr[3]), .ZN(n1899) );
  AOI211_X1 U1963 ( .C1(fmem_addr[3]), .C2(fmem_data[2]), .A(n1899), .B(n1845), 
        .ZN(n2518) );
  AOI22_X1 U1964 ( .A1(n1847), .A2(\xmem_inst/mem[24][10] ), .B1(n1846), .B2(
        \xmem_inst/mem[25][10] ), .ZN(n1857) );
  AOI22_X1 U1965 ( .A1(n1849), .A2(\xmem_inst/mem[0][10] ), .B1(n1848), .B2(
        \xmem_inst/mem[8][10] ), .ZN(n1856) );
  AOI22_X1 U1966 ( .A1(n1851), .A2(\xmem_inst/mem[16][10] ), .B1(n1850), .B2(
        \xmem_inst/mem[1][10] ), .ZN(n1855) );
  AOI22_X1 U1967 ( .A1(n1853), .A2(\xmem_inst/mem[9][10] ), .B1(n1852), .B2(
        \xmem_inst/mem[17][10] ), .ZN(n1854) );
  NAND4_X1 U1968 ( .A1(n1857), .A2(n1856), .A3(n1855), .A4(n1854), .ZN(n1882)
         );
  AOI22_X1 U1969 ( .A1(n1859), .A2(\xmem_inst/mem[26][10] ), .B1(n1858), .B2(
        \xmem_inst/mem[10][10] ), .ZN(n1869) );
  AOI22_X1 U1970 ( .A1(n1861), .A2(\xmem_inst/mem[2][10] ), .B1(n1860), .B2(
        \xmem_inst/mem[27][10] ), .ZN(n1868) );
  AOI22_X1 U1971 ( .A1(n1863), .A2(\xmem_inst/mem[18][10] ), .B1(n1862), .B2(
        \xmem_inst/mem[3][10] ), .ZN(n1867) );
  AOI22_X1 U1972 ( .A1(n1865), .A2(\xmem_inst/mem[11][10] ), .B1(n1864), .B2(
        \xmem_inst/mem[19][10] ), .ZN(n1866) );
  NAND4_X1 U1973 ( .A1(n1869), .A2(n1868), .A3(n1867), .A4(n1866), .ZN(n1881)
         );
  AOI22_X1 U1974 ( .A1(n1871), .A2(\xmem_inst/mem[28][10] ), .B1(n1870), .B2(
        \xmem_inst/mem[29][10] ), .ZN(n1879) );
  AOI22_X1 U1975 ( .A1(n1873), .A2(\xmem_inst/mem[4][10] ), .B1(n1872), .B2(
        \xmem_inst/mem[12][10] ), .ZN(n1878) );
  AOI22_X1 U1976 ( .A1(n2151), .A2(\xmem_inst/mem[14][10] ), .B1(n2043), .B2(
        \xmem_inst/mem[6][10] ), .ZN(n1877) );
  AOI22_X1 U1977 ( .A1(n1875), .A2(\xmem_inst/mem[20][10] ), .B1(n1874), .B2(
        \xmem_inst/mem[21][10] ), .ZN(n1876) );
  NAND4_X1 U1978 ( .A1(n1879), .A2(n1878), .A3(n1877), .A4(n1876), .ZN(n1880)
         );
  NOR3_X1 U1979 ( .A1(n1882), .A2(n1881), .A3(n1880), .ZN(n1889) );
  AOI22_X1 U1980 ( .A1(n1884), .A2(\xmem_inst/mem[5][10] ), .B1(n1883), .B2(
        \xmem_inst/mem[13][10] ), .ZN(n1888) );
  AOI22_X1 U1981 ( .A1(n1885), .A2(\xmem_inst/mem[15][10] ), .B1(n2275), .B2(
        \xmem_inst/mem[23][10] ), .ZN(n1887) );
  AOI22_X1 U1982 ( .A1(n2261), .A2(\xmem_inst/mem[22][10] ), .B1(n2057), .B2(
        \xmem_inst/mem[7][10] ), .ZN(n1886) );
  NAND4_X1 U1983 ( .A1(n1889), .A2(n1888), .A3(n1887), .A4(n1886), .ZN(
        \xmem_inst/N16 ) );
  NOR2_X1 U1984 ( .A1(n1944), .A2(n2379), .ZN(\ctrl_conv_output_inst/N74 ) );
  INV_X1 U1985 ( .A(\ctrl_conv_output_inst/N74 ), .ZN(n2380) );
  NOR3_X1 U1986 ( .A1(n2380), .A2(conv_done), .A3(
        \ctrl_conv_output_inst/m_pre_pre_valid_y ), .ZN(n1898) );
  INV_X1 U1987 ( .A(n1898), .ZN(n1892) );
  AOI21_X1 U1988 ( .B1(fmem_addr[3]), .B2(n1890), .A(n1892), .ZN(n1897) );
  INV_X1 U1989 ( .A(n1897), .ZN(n1895) );
  NAND2_X1 U1990 ( .A1(n1898), .A2(n2496), .ZN(n2374) );
  NOR2_X1 U1991 ( .A1(n1945), .A2(n1944), .ZN(n1891) );
  NOR2_X1 U1992 ( .A1(reset), .A2(conv_done), .ZN(n1939) );
  INV_X1 U1993 ( .A(n1939), .ZN(n1943) );
  NOR2_X1 U1994 ( .A1(n1891), .A2(n1943), .ZN(n1941) );
  NAND2_X1 U1995 ( .A1(n1941), .A2(n1892), .ZN(n2375) );
  NAND2_X1 U1996 ( .A1(n2374), .A2(n2375), .ZN(n1896) );
  INV_X1 U1997 ( .A(n1896), .ZN(n1893) );
  OAI22_X1 U1998 ( .A1(n1895), .A2(n1894), .B1(n1893), .B2(n2491), .ZN(n815)
         );
  NAND2_X1 U1999 ( .A1(n1897), .A2(n2489), .ZN(n2377) );
  AOI21_X1 U2000 ( .B1(n1897), .B2(n2491), .A(n1896), .ZN(n2378) );
  AND2_X1 U2001 ( .A1(n2377), .A2(n2378), .ZN(n1901) );
  NAND3_X1 U2002 ( .A1(fmem_addr[1]), .A2(n1899), .A3(n1898), .ZN(n1900) );
  OAI21_X1 U2003 ( .B1(n1901), .B2(n2498), .A(n1900), .ZN(n813) );
  NOR2_X1 U2004 ( .A1(\ctrl_conv_output_inst/m_pre_valid_y ), .A2(n2490), .ZN(
        n1925) );
  NAND2_X1 U2005 ( .A1(n1939), .A2(n1925), .ZN(n1928) );
  NAND2_X1 U2006 ( .A1(\ctrl_conv_output_inst/cnt_conv [1]), .A2(
        \ctrl_conv_output_inst/cnt_conv [0]), .ZN(n1924) );
  NOR2_X1 U2007 ( .A1(n1928), .A2(n1924), .ZN(n1904) );
  INV_X1 U2008 ( .A(n1928), .ZN(n1931) );
  AOI21_X1 U2009 ( .B1(\ctrl_conv_output_inst/cnt_conv [0]), .B2(n1925), .A(
        n1943), .ZN(n1930) );
  AOI21_X1 U2010 ( .B1(n1931), .B2(n2497), .A(n1930), .ZN(n1902) );
  INV_X1 U2011 ( .A(n1902), .ZN(n1903) );
  MUX2_X1 U2012 ( .A(n1904), .B(n1903), .S(\ctrl_conv_output_inst/cnt_conv [2]), .Z(n1155) );
  OR2_X1 U2013 ( .A1(n1906), .A2(n1177), .ZN(n1908) );
  NAND2_X1 U2014 ( .A1(n1906), .A2(n1177), .ZN(n1907) );
  NAND2_X1 U2015 ( .A1(n1908), .A2(n1907), .ZN(n1909) );
  XOR2_X1 U2016 ( .A(n1162), .B(n1909), .Z(n1918) );
  NAND2_X1 U2017 ( .A1(n1911), .A2(n1912), .ZN(n1917) );
  AOI21_X1 U2018 ( .B1(n1915), .B2(n1914), .A(n1244), .ZN(n1916) );
  OAI21_X1 U2019 ( .B1(n1917), .B2(n1918), .A(n1916), .ZN(n1919) );
  OAI21_X1 U2020 ( .B1(n2516), .B2(n1920), .A(n1919), .ZN(n795) );
  NAND4_X1 U2021 ( .A1(\ctrl_conv_output_inst/cnt_conv [1]), .A2(
        \ctrl_conv_output_inst/cnt_conv [4]), .A3(n2407), .A4(n2492), .ZN(
        n1921) );
  NOR4_X1 U2022 ( .A1(\ctrl_conv_output_inst/cnt_conv [3]), .A2(n2501), .A3(
        n1945), .A4(n1921), .ZN(\ctrl_conv_output_inst/N77 ) );
  AND2_X1 U2023 ( .A1(n2488), .A2(\mac_unit_inst/adder_reg [0]), .ZN(
        m_data_out_y[0]) );
  AND2_X1 U2024 ( .A1(n2488), .A2(\mac_unit_inst/adder_reg [1]), .ZN(
        m_data_out_y[1]) );
  AND2_X1 U2025 ( .A1(n2488), .A2(n2480), .ZN(m_data_out_y[2]) );
  AND2_X1 U2026 ( .A1(n2488), .A2(\mac_unit_inst/adder_reg [3]), .ZN(
        m_data_out_y[3]) );
  AND2_X1 U2027 ( .A1(n2488), .A2(\mac_unit_inst/adder_reg [4]), .ZN(
        m_data_out_y[4]) );
  AND2_X1 U2028 ( .A1(n2488), .A2(\mac_unit_inst/adder_reg [5]), .ZN(
        m_data_out_y[5]) );
  AND2_X1 U2029 ( .A1(n2488), .A2(\mac_unit_inst/adder_reg [6]), .ZN(
        m_data_out_y[6]) );
  AND2_X1 U2030 ( .A1(n2488), .A2(\mac_unit_inst/adder_reg [7]), .ZN(
        m_data_out_y[7]) );
  AND2_X1 U2031 ( .A1(n2488), .A2(\mac_unit_inst/adder_reg [8]), .ZN(
        m_data_out_y[8]) );
  AND2_X1 U2032 ( .A1(n2488), .A2(\mac_unit_inst/adder_reg [9]), .ZN(
        m_data_out_y[9]) );
  NOR2_X1 U2034 ( .A1(s_ready_x), .A2(reset), .ZN(N29) );
  NAND4_X1 U2035 ( .A1(n1940), .A2(fmem_addr[3]), .A3(n2490), .A4(n2407), .ZN(
        n1922) );
  OAI22_X1 U2036 ( .A1(n2490), .A2(n2379), .B1(n1923), .B2(n1922), .ZN(n1159)
         );
  NOR2_X1 U2037 ( .A1(n2501), .A2(n1924), .ZN(n1934) );
  NAND3_X1 U2038 ( .A1(\ctrl_conv_output_inst/cnt_conv [3]), .A2(n1931), .A3(
        n1934), .ZN(n1927) );
  AOI21_X1 U2039 ( .B1(n1925), .B2(n1934), .A(n1943), .ZN(n1936) );
  NOR2_X1 U2040 ( .A1(\ctrl_conv_output_inst/cnt_conv [3]), .A2(n1928), .ZN(
        n1935) );
  OAI21_X1 U2041 ( .B1(n1936), .B2(n1935), .A(
        \ctrl_conv_output_inst/cnt_conv [4]), .ZN(n1926) );
  OAI21_X1 U2042 ( .B1(\ctrl_conv_output_inst/cnt_conv [4]), .B2(n1927), .A(
        n1926), .ZN(n1158) );
  OAI21_X1 U2043 ( .B1(\ctrl_conv_output_inst/m_pre_valid_y ), .B2(n2490), .A(
        n1939), .ZN(n1929) );
  AOI22_X1 U2044 ( .A1(\ctrl_conv_output_inst/cnt_conv [0]), .A2(n1929), .B1(
        n1928), .B2(n2492), .ZN(n1157) );
  INV_X1 U2045 ( .A(n1930), .ZN(n1933) );
  NAND2_X1 U2046 ( .A1(n1931), .A2(n2497), .ZN(n1932) );
  OAI22_X1 U2047 ( .A1(n1933), .A2(n2497), .B1(n2492), .B2(n1932), .ZN(n1156)
         );
  AOI22_X1 U2048 ( .A1(\ctrl_conv_output_inst/cnt_conv [3]), .A2(n1936), .B1(
        n1935), .B2(n1934), .ZN(n2519) );
  NAND2_X1 U2049 ( .A1(m_valid_y), .A2(n2407), .ZN(n1937) );
  OAI22_X1 U2050 ( .A1(m_ready_y), .A2(n1937), .B1(n2503), .B2(n2380), .ZN(
        n1153) );
  NOR2_X2 U2051 ( .A1(n2247), .A2(n2347), .ZN(n2371) );
  OAI21_X1 U2052 ( .B1(n2371), .B2(n2511), .A(n1939), .ZN(n1152) );
  NAND3_X1 U2053 ( .A1(n1940), .A2(n1945), .A3(n2490), .ZN(n1942) );
  NAND3_X1 U2054 ( .A1(n1941), .A2(n2166), .A3(n1942), .ZN(n1954) );
  AOI211_X1 U2055 ( .C1(n1942), .C2(n2166), .A(n2371), .B(n1943), .ZN(n1953)
         );
  NAND2_X1 U2056 ( .A1(n1953), .A2(n2493), .ZN(n1947) );
  NOR3_X1 U2057 ( .A1(n1945), .A2(n1944), .A3(n1943), .ZN(n1958) );
  NAND2_X1 U2058 ( .A1(n1958), .A2(\ctrl_conv_output_inst/cnt_conv [0]), .ZN(
        n1946) );
  OAI211_X1 U2059 ( .C1(n2493), .C2(n1954), .A(n1947), .B(n1946), .ZN(n1151)
         );
  NAND2_X1 U2060 ( .A1(n1953), .A2(xmem_addr[0]), .ZN(n1949) );
  NAND2_X1 U2061 ( .A1(n1954), .A2(n1947), .ZN(n1950) );
  AOI22_X1 U2062 ( .A1(xmem_addr[1]), .A2(n1950), .B1(n1958), .B2(
        \ctrl_conv_output_inst/cnt_conv [1]), .ZN(n1948) );
  OAI21_X1 U2063 ( .B1(n1949), .B2(xmem_addr[1]), .A(n1948), .ZN(n1150) );
  INV_X1 U2064 ( .A(n1953), .ZN(n1962) );
  AOI22_X1 U2065 ( .A1(xmem_addr[2]), .A2(n1950), .B1(n1958), .B2(
        \ctrl_conv_output_inst/cnt_conv [2]), .ZN(n1951) );
  OAI221_X1 U2066 ( .B1(n1962), .B2(n1952), .C1(n1962), .C2(n2332), .A(n1951), 
        .ZN(n1149) );
  NAND3_X1 U2067 ( .A1(n2495), .A2(n1955), .A3(n1953), .ZN(n1957) );
  OAI21_X1 U2068 ( .B1(n1955), .B2(n1962), .A(n1954), .ZN(n1959) );
  AOI22_X1 U2069 ( .A1(xmem_addr[3]), .A2(n1959), .B1(n1958), .B2(
        \ctrl_conv_output_inst/cnt_conv [3]), .ZN(n1956) );
  NAND2_X1 U2070 ( .A1(n1957), .A2(n1956), .ZN(n1148) );
  AOI22_X1 U2071 ( .A1(xmem_addr[4]), .A2(n1959), .B1(n1958), .B2(
        \ctrl_conv_output_inst/cnt_conv [4]), .ZN(n1960) );
  OAI221_X1 U2072 ( .B1(n1962), .B2(n1961), .C1(n1962), .C2(n2165), .A(n1960), 
        .ZN(n1147) );
  NAND2_X1 U2073 ( .A1(n2276), .A2(n1963), .ZN(n2029) );
  NOR2_X1 U2074 ( .A1(n2290), .A2(n2029), .ZN(n1974) );
  INV_X1 U2075 ( .A(n1974), .ZN(n1975) );
  OAI22_X1 U2076 ( .A1(n1975), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[0][0] ), 
        .B2(n1974), .ZN(n1964) );
  INV_X1 U2077 ( .A(n1964), .ZN(n1146) );
  OAI22_X1 U2078 ( .A1(n1975), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[0][1] ), 
        .B2(n1974), .ZN(n1965) );
  INV_X1 U2079 ( .A(n1965), .ZN(n1145) );
  OAI22_X1 U2080 ( .A1(n1975), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[0][2] ), 
        .B2(n1974), .ZN(n1966) );
  INV_X1 U2081 ( .A(n1966), .ZN(n1144) );
  OAI22_X1 U2082 ( .A1(n1975), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[0][3] ), 
        .B2(n1974), .ZN(n1967) );
  INV_X1 U2083 ( .A(n1967), .ZN(n1143) );
  OAI22_X1 U2084 ( .A1(n1975), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[0][4] ), 
        .B2(n1974), .ZN(n1968) );
  INV_X1 U2085 ( .A(n1968), .ZN(n1142) );
  OAI22_X1 U2086 ( .A1(n1975), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[0][5] ), 
        .B2(n1974), .ZN(n1969) );
  INV_X1 U2087 ( .A(n1969), .ZN(n1141) );
  OAI22_X1 U2088 ( .A1(n1975), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[0][6] ), 
        .B2(n1974), .ZN(n1970) );
  INV_X1 U2089 ( .A(n1970), .ZN(n1140) );
  OAI22_X1 U2090 ( .A1(n1975), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[0][7] ), 
        .B2(n1974), .ZN(n1971) );
  INV_X1 U2091 ( .A(n1971), .ZN(n1139) );
  OAI22_X1 U2092 ( .A1(n1975), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[0][8] ), 
        .B2(n1974), .ZN(n1972) );
  INV_X1 U2093 ( .A(n1972), .ZN(n1138) );
  OAI22_X1 U2094 ( .A1(n1975), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[0][9] ), 
        .B2(n1974), .ZN(n1973) );
  INV_X1 U2095 ( .A(n1973), .ZN(n1137) );
  OAI22_X1 U2096 ( .A1(n1975), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[0][10] ), .B2(n1974), .ZN(n1976) );
  INV_X1 U2097 ( .A(n1976), .ZN(n1136) );
  NOR2_X1 U2098 ( .A1(n2304), .A2(n2029), .ZN(n1987) );
  INV_X1 U2099 ( .A(n1987), .ZN(n1988) );
  OAI22_X1 U2100 ( .A1(n1988), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[1][0] ), 
        .B2(n1987), .ZN(n1977) );
  INV_X1 U2101 ( .A(n1977), .ZN(n1135) );
  OAI22_X1 U2102 ( .A1(n1988), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[1][1] ), 
        .B2(n1987), .ZN(n1978) );
  INV_X1 U2103 ( .A(n1978), .ZN(n1134) );
  OAI22_X1 U2104 ( .A1(n1988), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[1][2] ), 
        .B2(n1987), .ZN(n1979) );
  INV_X1 U2105 ( .A(n1979), .ZN(n1133) );
  OAI22_X1 U2106 ( .A1(n1988), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[1][3] ), 
        .B2(n1987), .ZN(n1980) );
  INV_X1 U2107 ( .A(n1980), .ZN(n1132) );
  OAI22_X1 U2108 ( .A1(n1988), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[1][4] ), 
        .B2(n1987), .ZN(n1981) );
  INV_X1 U2109 ( .A(n1981), .ZN(n1131) );
  OAI22_X1 U2110 ( .A1(n1988), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[1][5] ), 
        .B2(n1987), .ZN(n1982) );
  INV_X1 U2111 ( .A(n1982), .ZN(n1130) );
  OAI22_X1 U2112 ( .A1(n1988), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[1][6] ), 
        .B2(n1987), .ZN(n1983) );
  INV_X1 U2113 ( .A(n1983), .ZN(n1129) );
  OAI22_X1 U2114 ( .A1(n1988), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[1][7] ), 
        .B2(n1987), .ZN(n1984) );
  INV_X1 U2115 ( .A(n1984), .ZN(n1128) );
  OAI22_X1 U2116 ( .A1(n1988), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[1][8] ), 
        .B2(n1987), .ZN(n1985) );
  INV_X1 U2117 ( .A(n1985), .ZN(n1127) );
  OAI22_X1 U2118 ( .A1(n1988), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[1][9] ), 
        .B2(n1987), .ZN(n1986) );
  INV_X1 U2119 ( .A(n1986), .ZN(n1126) );
  OAI22_X1 U2120 ( .A1(n1988), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[1][10] ), .B2(n1987), .ZN(n1989) );
  INV_X1 U2121 ( .A(n1989), .ZN(n1125) );
  NOR2_X1 U2122 ( .A1(n2318), .A2(n2029), .ZN(n2000) );
  INV_X1 U2123 ( .A(n2000), .ZN(n2001) );
  OAI22_X1 U2124 ( .A1(n2001), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[2][0] ), 
        .B2(n2000), .ZN(n1990) );
  INV_X1 U2125 ( .A(n1990), .ZN(n1124) );
  OAI22_X1 U2126 ( .A1(n2001), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[2][1] ), 
        .B2(n2000), .ZN(n1991) );
  INV_X1 U2127 ( .A(n1991), .ZN(n1123) );
  OAI22_X1 U2128 ( .A1(n2001), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[2][2] ), 
        .B2(n2000), .ZN(n1992) );
  INV_X1 U2129 ( .A(n1992), .ZN(n1122) );
  OAI22_X1 U2130 ( .A1(n2001), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[2][3] ), 
        .B2(n2000), .ZN(n1993) );
  INV_X1 U2131 ( .A(n1993), .ZN(n1121) );
  OAI22_X1 U2132 ( .A1(n2001), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[2][4] ), 
        .B2(n2000), .ZN(n1994) );
  INV_X1 U2133 ( .A(n1994), .ZN(n1120) );
  OAI22_X1 U2134 ( .A1(n2001), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[2][5] ), 
        .B2(n2000), .ZN(n1995) );
  INV_X1 U2135 ( .A(n1995), .ZN(n1119) );
  OAI22_X1 U2136 ( .A1(n2001), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[2][6] ), 
        .B2(n2000), .ZN(n1996) );
  INV_X1 U2137 ( .A(n1996), .ZN(n1118) );
  OAI22_X1 U2138 ( .A1(n2001), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[2][7] ), 
        .B2(n2000), .ZN(n1997) );
  INV_X1 U2139 ( .A(n1997), .ZN(n1117) );
  OAI22_X1 U2140 ( .A1(n2001), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[2][8] ), 
        .B2(n2000), .ZN(n1998) );
  INV_X1 U2141 ( .A(n1998), .ZN(n1116) );
  OAI22_X1 U2142 ( .A1(n2001), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[2][9] ), 
        .B2(n2000), .ZN(n1999) );
  INV_X1 U2143 ( .A(n1999), .ZN(n1115) );
  OAI22_X1 U2144 ( .A1(n2001), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[2][10] ), .B2(n2000), .ZN(n2002) );
  INV_X1 U2145 ( .A(n2002), .ZN(n1114) );
  NOR2_X1 U2146 ( .A1(n2332), .A2(n2029), .ZN(n2013) );
  INV_X1 U2147 ( .A(n2013), .ZN(n2014) );
  OAI22_X1 U2148 ( .A1(n2014), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[3][0] ), 
        .B2(n2013), .ZN(n2003) );
  INV_X1 U2149 ( .A(n2003), .ZN(n1113) );
  OAI22_X1 U2150 ( .A1(n2014), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[3][1] ), 
        .B2(n2013), .ZN(n2004) );
  INV_X1 U2151 ( .A(n2004), .ZN(n1112) );
  OAI22_X1 U2152 ( .A1(n2014), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[3][2] ), 
        .B2(n2013), .ZN(n2005) );
  INV_X1 U2153 ( .A(n2005), .ZN(n1111) );
  OAI22_X1 U2154 ( .A1(n2014), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[3][3] ), 
        .B2(n2013), .ZN(n2006) );
  INV_X1 U2155 ( .A(n2006), .ZN(n1110) );
  OAI22_X1 U2156 ( .A1(n2014), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[3][4] ), 
        .B2(n2013), .ZN(n2007) );
  INV_X1 U2157 ( .A(n2007), .ZN(n1109) );
  OAI22_X1 U2158 ( .A1(n2014), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[3][5] ), 
        .B2(n2013), .ZN(n2008) );
  INV_X1 U2159 ( .A(n2008), .ZN(n1108) );
  OAI22_X1 U2160 ( .A1(n2014), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[3][6] ), 
        .B2(n2013), .ZN(n2009) );
  INV_X1 U2161 ( .A(n2009), .ZN(n1107) );
  OAI22_X1 U2162 ( .A1(n2014), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[3][7] ), 
        .B2(n2013), .ZN(n2010) );
  INV_X1 U2163 ( .A(n2010), .ZN(n1106) );
  OAI22_X1 U2164 ( .A1(n2014), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[3][8] ), 
        .B2(n2013), .ZN(n2011) );
  INV_X1 U2165 ( .A(n2011), .ZN(n1105) );
  OAI22_X1 U2166 ( .A1(n2014), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[3][9] ), 
        .B2(n2013), .ZN(n2012) );
  INV_X1 U2167 ( .A(n2012), .ZN(n1104) );
  OAI22_X1 U2168 ( .A1(n2014), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[3][10] ), .B2(n2013), .ZN(n2015) );
  INV_X1 U2169 ( .A(n2015), .ZN(n1103) );
  NOR2_X1 U2170 ( .A1(n2346), .A2(n2029), .ZN(n2026) );
  INV_X1 U2171 ( .A(n2026), .ZN(n2027) );
  OAI22_X1 U2172 ( .A1(n2027), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[4][0] ), 
        .B2(n2026), .ZN(n2016) );
  INV_X1 U2173 ( .A(n2016), .ZN(n1102) );
  OAI22_X1 U2174 ( .A1(n2027), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[4][1] ), 
        .B2(n2026), .ZN(n2017) );
  INV_X1 U2175 ( .A(n2017), .ZN(n1101) );
  OAI22_X1 U2176 ( .A1(n2027), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[4][2] ), 
        .B2(n2026), .ZN(n2018) );
  INV_X1 U2177 ( .A(n2018), .ZN(n1100) );
  OAI22_X1 U2178 ( .A1(n2027), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[4][3] ), 
        .B2(n2026), .ZN(n2019) );
  INV_X1 U2179 ( .A(n2019), .ZN(n1099) );
  OAI22_X1 U2180 ( .A1(n2027), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[4][4] ), 
        .B2(n2026), .ZN(n2020) );
  INV_X1 U2181 ( .A(n2020), .ZN(n1098) );
  OAI22_X1 U2182 ( .A1(n2027), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[4][5] ), 
        .B2(n2026), .ZN(n2021) );
  INV_X1 U2183 ( .A(n2021), .ZN(n1097) );
  OAI22_X1 U2184 ( .A1(n2027), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[4][6] ), 
        .B2(n2026), .ZN(n2022) );
  INV_X1 U2185 ( .A(n2022), .ZN(n1096) );
  OAI22_X1 U2186 ( .A1(n2027), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[4][7] ), 
        .B2(n2026), .ZN(n2023) );
  INV_X1 U2187 ( .A(n2023), .ZN(n1095) );
  OAI22_X1 U2188 ( .A1(n2027), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[4][8] ), 
        .B2(n2026), .ZN(n2024) );
  INV_X1 U2189 ( .A(n2024), .ZN(n1094) );
  OAI22_X1 U2190 ( .A1(n2027), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[4][9] ), 
        .B2(n2026), .ZN(n2025) );
  INV_X1 U2191 ( .A(n2025), .ZN(n1093) );
  OAI22_X1 U2192 ( .A1(n2027), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[4][10] ), .B2(n2026), .ZN(n2028) );
  INV_X1 U2193 ( .A(n2028), .ZN(n1092) );
  NOR2_X1 U2194 ( .A1(n2247), .A2(n2029), .ZN(n2040) );
  INV_X1 U2195 ( .A(n2040), .ZN(n2041) );
  OAI22_X1 U2196 ( .A1(n2041), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[5][0] ), 
        .B2(n2040), .ZN(n2030) );
  INV_X1 U2197 ( .A(n2030), .ZN(n1091) );
  OAI22_X1 U2198 ( .A1(n2041), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[5][1] ), 
        .B2(n2040), .ZN(n2031) );
  INV_X1 U2199 ( .A(n2031), .ZN(n1090) );
  OAI22_X1 U2200 ( .A1(n2041), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[5][2] ), 
        .B2(n2040), .ZN(n2032) );
  INV_X1 U2201 ( .A(n2032), .ZN(n1089) );
  OAI22_X1 U2202 ( .A1(n2041), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[5][3] ), 
        .B2(n2040), .ZN(n2033) );
  INV_X1 U2203 ( .A(n2033), .ZN(n1088) );
  OAI22_X1 U2204 ( .A1(n2041), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[5][4] ), 
        .B2(n2040), .ZN(n2034) );
  INV_X1 U2205 ( .A(n2034), .ZN(n1087) );
  OAI22_X1 U2206 ( .A1(n2041), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[5][5] ), 
        .B2(n2040), .ZN(n2035) );
  INV_X1 U2207 ( .A(n2035), .ZN(n1086) );
  OAI22_X1 U2208 ( .A1(n2041), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[5][6] ), 
        .B2(n2040), .ZN(n2036) );
  INV_X1 U2209 ( .A(n2036), .ZN(n1085) );
  OAI22_X1 U2210 ( .A1(n2041), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[5][7] ), 
        .B2(n2040), .ZN(n2037) );
  INV_X1 U2211 ( .A(n2037), .ZN(n1084) );
  OAI22_X1 U2212 ( .A1(n2041), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[5][8] ), 
        .B2(n2040), .ZN(n2038) );
  INV_X1 U2213 ( .A(n2038), .ZN(n1083) );
  OAI22_X1 U2214 ( .A1(n2041), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[5][9] ), 
        .B2(n2040), .ZN(n2039) );
  INV_X1 U2215 ( .A(n2039), .ZN(n1082) );
  OAI22_X1 U2216 ( .A1(n2041), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[5][10] ), .B2(n2040), .ZN(n2042) );
  INV_X1 U2217 ( .A(n2042), .ZN(n1081) );
  NAND2_X1 U2218 ( .A1(n2276), .A2(n2043), .ZN(n2055) );
  OAI22_X1 U2219 ( .A1(n2055), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[6][0] ), 
        .B2(n2054), .ZN(n2044) );
  INV_X1 U2220 ( .A(n2044), .ZN(n1080) );
  OAI22_X1 U2221 ( .A1(n2055), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[6][1] ), 
        .B2(n2054), .ZN(n2045) );
  INV_X1 U2222 ( .A(n2045), .ZN(n1079) );
  OAI22_X1 U2223 ( .A1(n2055), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[6][2] ), 
        .B2(n2054), .ZN(n2046) );
  INV_X1 U2224 ( .A(n2046), .ZN(n1078) );
  OAI22_X1 U2225 ( .A1(n2055), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[6][3] ), 
        .B2(n2054), .ZN(n2047) );
  INV_X1 U2226 ( .A(n2047), .ZN(n1077) );
  OAI22_X1 U2227 ( .A1(n2055), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[6][4] ), 
        .B2(n2054), .ZN(n2048) );
  INV_X1 U2228 ( .A(n2048), .ZN(n1076) );
  OAI22_X1 U2229 ( .A1(n2055), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[6][5] ), 
        .B2(n2054), .ZN(n2049) );
  INV_X1 U2230 ( .A(n2049), .ZN(n1075) );
  OAI22_X1 U2231 ( .A1(n2055), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[6][6] ), 
        .B2(n2054), .ZN(n2050) );
  INV_X1 U2232 ( .A(n2050), .ZN(n1074) );
  OAI22_X1 U2233 ( .A1(n2055), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[6][7] ), 
        .B2(n2054), .ZN(n2051) );
  INV_X1 U2234 ( .A(n2051), .ZN(n1073) );
  OAI22_X1 U2235 ( .A1(n2055), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[6][8] ), 
        .B2(n2054), .ZN(n2052) );
  INV_X1 U2236 ( .A(n2052), .ZN(n1072) );
  OAI22_X1 U2237 ( .A1(n2055), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[6][9] ), 
        .B2(n2054), .ZN(n2053) );
  INV_X1 U2238 ( .A(n2053), .ZN(n1071) );
  OAI22_X1 U2239 ( .A1(n2055), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[6][10] ), .B2(n2054), .ZN(n2056) );
  INV_X1 U2240 ( .A(n2056), .ZN(n1070) );
  NAND2_X1 U2241 ( .A1(n2276), .A2(n2057), .ZN(n2069) );
  OAI22_X1 U2242 ( .A1(n2069), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[7][0] ), 
        .B2(n2068), .ZN(n2058) );
  INV_X1 U2243 ( .A(n2058), .ZN(n1069) );
  OAI22_X1 U2244 ( .A1(n2069), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[7][1] ), 
        .B2(n2068), .ZN(n2059) );
  INV_X1 U2245 ( .A(n2059), .ZN(n1068) );
  OAI22_X1 U2246 ( .A1(n2069), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[7][2] ), 
        .B2(n2068), .ZN(n2060) );
  INV_X1 U2247 ( .A(n2060), .ZN(n1067) );
  OAI22_X1 U2248 ( .A1(n2069), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[7][3] ), 
        .B2(n2068), .ZN(n2061) );
  INV_X1 U2249 ( .A(n2061), .ZN(n1066) );
  OAI22_X1 U2250 ( .A1(n2069), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[7][4] ), 
        .B2(n2068), .ZN(n2062) );
  INV_X1 U2251 ( .A(n2062), .ZN(n1065) );
  OAI22_X1 U2252 ( .A1(n2069), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[7][5] ), 
        .B2(n2068), .ZN(n2063) );
  INV_X1 U2253 ( .A(n2063), .ZN(n1064) );
  OAI22_X1 U2254 ( .A1(n2069), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[7][6] ), 
        .B2(n2068), .ZN(n2064) );
  INV_X1 U2255 ( .A(n2064), .ZN(n1063) );
  OAI22_X1 U2256 ( .A1(n2069), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[7][7] ), 
        .B2(n2068), .ZN(n2065) );
  INV_X1 U2257 ( .A(n2065), .ZN(n1062) );
  OAI22_X1 U2258 ( .A1(n2069), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[7][8] ), 
        .B2(n2068), .ZN(n2066) );
  INV_X1 U2259 ( .A(n2066), .ZN(n1061) );
  OAI22_X1 U2260 ( .A1(n2069), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[7][9] ), 
        .B2(n2068), .ZN(n2067) );
  INV_X1 U2261 ( .A(n2067), .ZN(n1060) );
  OAI22_X1 U2262 ( .A1(n2069), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[7][10] ), .B2(n2068), .ZN(n2070) );
  INV_X1 U2263 ( .A(n2070), .ZN(n1059) );
  NAND2_X1 U2264 ( .A1(n2276), .A2(n2071), .ZN(n2137) );
  NOR2_X1 U2265 ( .A1(n2290), .A2(n2137), .ZN(n2082) );
  INV_X1 U2266 ( .A(n2082), .ZN(n2083) );
  OAI22_X1 U2267 ( .A1(n2083), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[8][0] ), 
        .B2(n2082), .ZN(n2072) );
  INV_X1 U2268 ( .A(n2072), .ZN(n1058) );
  OAI22_X1 U2269 ( .A1(n2083), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[8][1] ), 
        .B2(n2082), .ZN(n2073) );
  INV_X1 U2270 ( .A(n2073), .ZN(n1057) );
  OAI22_X1 U2271 ( .A1(n2083), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[8][2] ), 
        .B2(n2082), .ZN(n2074) );
  INV_X1 U2272 ( .A(n2074), .ZN(n1056) );
  OAI22_X1 U2273 ( .A1(n2083), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[8][3] ), 
        .B2(n2082), .ZN(n2075) );
  INV_X1 U2274 ( .A(n2075), .ZN(n1055) );
  OAI22_X1 U2275 ( .A1(n2083), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[8][4] ), 
        .B2(n2082), .ZN(n2076) );
  INV_X1 U2276 ( .A(n2076), .ZN(n1054) );
  OAI22_X1 U2277 ( .A1(n2083), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[8][5] ), 
        .B2(n2082), .ZN(n2077) );
  INV_X1 U2278 ( .A(n2077), .ZN(n1053) );
  OAI22_X1 U2279 ( .A1(n2083), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[8][6] ), 
        .B2(n2082), .ZN(n2078) );
  INV_X1 U2280 ( .A(n2078), .ZN(n1052) );
  OAI22_X1 U2281 ( .A1(n2083), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[8][7] ), 
        .B2(n2082), .ZN(n2079) );
  INV_X1 U2282 ( .A(n2079), .ZN(n1051) );
  OAI22_X1 U2283 ( .A1(n2083), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[8][8] ), 
        .B2(n2082), .ZN(n2080) );
  INV_X1 U2284 ( .A(n2080), .ZN(n1050) );
  OAI22_X1 U2285 ( .A1(n2083), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[8][9] ), 
        .B2(n2082), .ZN(n2081) );
  INV_X1 U2286 ( .A(n2081), .ZN(n1049) );
  OAI22_X1 U2287 ( .A1(n2083), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[8][10] ), .B2(n2082), .ZN(n2084) );
  INV_X1 U2288 ( .A(n2084), .ZN(n1048) );
  NOR2_X1 U2289 ( .A1(n2304), .A2(n2137), .ZN(n2095) );
  INV_X1 U2290 ( .A(n2095), .ZN(n2096) );
  OAI22_X1 U2291 ( .A1(n2096), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[9][0] ), 
        .B2(n2095), .ZN(n2085) );
  INV_X1 U2292 ( .A(n2085), .ZN(n1047) );
  OAI22_X1 U2293 ( .A1(n2096), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[9][1] ), 
        .B2(n2095), .ZN(n2086) );
  INV_X1 U2294 ( .A(n2086), .ZN(n1046) );
  OAI22_X1 U2295 ( .A1(n2096), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[9][2] ), 
        .B2(n2095), .ZN(n2087) );
  INV_X1 U2296 ( .A(n2087), .ZN(n1045) );
  OAI22_X1 U2297 ( .A1(n2096), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[9][3] ), 
        .B2(n2095), .ZN(n2088) );
  INV_X1 U2298 ( .A(n2088), .ZN(n1044) );
  OAI22_X1 U2299 ( .A1(n2096), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[9][4] ), 
        .B2(n2095), .ZN(n2089) );
  INV_X1 U2300 ( .A(n2089), .ZN(n1043) );
  OAI22_X1 U2301 ( .A1(n2096), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[9][5] ), 
        .B2(n2095), .ZN(n2090) );
  INV_X1 U2302 ( .A(n2090), .ZN(n1042) );
  OAI22_X1 U2303 ( .A1(n2096), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[9][6] ), 
        .B2(n2095), .ZN(n2091) );
  INV_X1 U2304 ( .A(n2091), .ZN(n1041) );
  OAI22_X1 U2305 ( .A1(n2096), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[9][7] ), 
        .B2(n2095), .ZN(n2092) );
  INV_X1 U2306 ( .A(n2092), .ZN(n1040) );
  OAI22_X1 U2307 ( .A1(n2096), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[9][8] ), 
        .B2(n2095), .ZN(n2093) );
  INV_X1 U2308 ( .A(n2093), .ZN(n1039) );
  OAI22_X1 U2309 ( .A1(n2096), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[9][9] ), 
        .B2(n2095), .ZN(n2094) );
  INV_X1 U2310 ( .A(n2094), .ZN(n1038) );
  OAI22_X1 U2311 ( .A1(n2096), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[9][10] ), .B2(n2095), .ZN(n2097) );
  INV_X1 U2312 ( .A(n2097), .ZN(n1037) );
  NOR2_X1 U2313 ( .A1(n2318), .A2(n2137), .ZN(n2108) );
  INV_X1 U2314 ( .A(n2108), .ZN(n2109) );
  OAI22_X1 U2315 ( .A1(n2109), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[10][0] ), .B2(n2108), .ZN(n2098) );
  INV_X1 U2316 ( .A(n2098), .ZN(n1036) );
  OAI22_X1 U2317 ( .A1(n2109), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[10][1] ), .B2(n2108), .ZN(n2099) );
  INV_X1 U2318 ( .A(n2099), .ZN(n1035) );
  OAI22_X1 U2319 ( .A1(n2109), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[10][2] ), .B2(n2108), .ZN(n2100) );
  INV_X1 U2320 ( .A(n2100), .ZN(n1034) );
  OAI22_X1 U2321 ( .A1(n2109), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[10][3] ), .B2(n2108), .ZN(n2101) );
  INV_X1 U2322 ( .A(n2101), .ZN(n1033) );
  OAI22_X1 U2323 ( .A1(n2109), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[10][4] ), .B2(n2108), .ZN(n2102) );
  INV_X1 U2324 ( .A(n2102), .ZN(n1032) );
  OAI22_X1 U2325 ( .A1(n2109), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[10][5] ), .B2(n2108), .ZN(n2103) );
  INV_X1 U2326 ( .A(n2103), .ZN(n1031) );
  OAI22_X1 U2327 ( .A1(n2109), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[10][6] ), .B2(n2108), .ZN(n2104) );
  INV_X1 U2328 ( .A(n2104), .ZN(n1030) );
  OAI22_X1 U2329 ( .A1(n2109), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[10][7] ), .B2(n2108), .ZN(n2105) );
  INV_X1 U2330 ( .A(n2105), .ZN(n1029) );
  OAI22_X1 U2331 ( .A1(n2109), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[10][8] ), .B2(n2108), .ZN(n2106) );
  INV_X1 U2332 ( .A(n2106), .ZN(n1028) );
  OAI22_X1 U2333 ( .A1(n2109), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[10][9] ), .B2(n2108), .ZN(n2107) );
  INV_X1 U2334 ( .A(n2107), .ZN(n1027) );
  OAI22_X1 U2335 ( .A1(n2109), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[10][10] ), .B2(n2108), .ZN(n2110) );
  INV_X1 U2336 ( .A(n2110), .ZN(n1026) );
  NOR2_X1 U2337 ( .A1(n2332), .A2(n2137), .ZN(n2121) );
  INV_X1 U2338 ( .A(n2121), .ZN(n2122) );
  OAI22_X1 U2339 ( .A1(n2122), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[11][0] ), .B2(n2121), .ZN(n2111) );
  INV_X1 U2340 ( .A(n2111), .ZN(n1025) );
  OAI22_X1 U2341 ( .A1(n2122), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[11][1] ), .B2(n2121), .ZN(n2112) );
  INV_X1 U2342 ( .A(n2112), .ZN(n1024) );
  OAI22_X1 U2343 ( .A1(n2122), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[11][2] ), .B2(n2121), .ZN(n2113) );
  INV_X1 U2344 ( .A(n2113), .ZN(n1023) );
  OAI22_X1 U2345 ( .A1(n2122), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[11][3] ), .B2(n2121), .ZN(n2114) );
  INV_X1 U2346 ( .A(n2114), .ZN(n1022) );
  OAI22_X1 U2347 ( .A1(n2122), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[11][4] ), .B2(n2121), .ZN(n2115) );
  INV_X1 U2348 ( .A(n2115), .ZN(n1021) );
  OAI22_X1 U2349 ( .A1(n2122), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[11][5] ), .B2(n2121), .ZN(n2116) );
  INV_X1 U2350 ( .A(n2116), .ZN(n1020) );
  OAI22_X1 U2351 ( .A1(n2122), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[11][6] ), .B2(n2121), .ZN(n2117) );
  INV_X1 U2352 ( .A(n2117), .ZN(n1019) );
  OAI22_X1 U2353 ( .A1(n2122), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[11][7] ), .B2(n2121), .ZN(n2118) );
  INV_X1 U2354 ( .A(n2118), .ZN(n1018) );
  OAI22_X1 U2355 ( .A1(n2122), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[11][8] ), .B2(n2121), .ZN(n2119) );
  INV_X1 U2356 ( .A(n2119), .ZN(n1017) );
  OAI22_X1 U2357 ( .A1(n2122), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[11][9] ), .B2(n2121), .ZN(n2120) );
  INV_X1 U2358 ( .A(n2120), .ZN(n1016) );
  OAI22_X1 U2359 ( .A1(n2122), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[11][10] ), .B2(n2121), .ZN(n2123) );
  INV_X1 U2360 ( .A(n2123), .ZN(n1015) );
  NOR2_X1 U2361 ( .A1(n2346), .A2(n2137), .ZN(n2134) );
  INV_X1 U2362 ( .A(n2134), .ZN(n2135) );
  OAI22_X1 U2363 ( .A1(n2135), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[12][0] ), .B2(n2134), .ZN(n2124) );
  INV_X1 U2364 ( .A(n2124), .ZN(n1014) );
  OAI22_X1 U2365 ( .A1(n2135), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[12][1] ), .B2(n2134), .ZN(n2125) );
  INV_X1 U2366 ( .A(n2125), .ZN(n1013) );
  OAI22_X1 U2367 ( .A1(n2135), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[12][2] ), .B2(n2134), .ZN(n2126) );
  INV_X1 U2368 ( .A(n2126), .ZN(n1012) );
  OAI22_X1 U2369 ( .A1(n2135), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[12][3] ), .B2(n2134), .ZN(n2127) );
  INV_X1 U2370 ( .A(n2127), .ZN(n1011) );
  OAI22_X1 U2371 ( .A1(n2135), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[12][4] ), .B2(n2134), .ZN(n2128) );
  INV_X1 U2372 ( .A(n2128), .ZN(n1010) );
  OAI22_X1 U2373 ( .A1(n2135), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[12][5] ), .B2(n2134), .ZN(n2129) );
  INV_X1 U2374 ( .A(n2129), .ZN(n1009) );
  OAI22_X1 U2375 ( .A1(n2135), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[12][6] ), .B2(n2134), .ZN(n2130) );
  INV_X1 U2376 ( .A(n2130), .ZN(n1008) );
  OAI22_X1 U2377 ( .A1(n2135), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[12][7] ), .B2(n2134), .ZN(n2131) );
  INV_X1 U2378 ( .A(n2131), .ZN(n1007) );
  OAI22_X1 U2379 ( .A1(n2135), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[12][8] ), .B2(n2134), .ZN(n2132) );
  INV_X1 U2380 ( .A(n2132), .ZN(n1006) );
  OAI22_X1 U2381 ( .A1(n2135), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[12][9] ), .B2(n2134), .ZN(n2133) );
  INV_X1 U2382 ( .A(n2133), .ZN(n1005) );
  OAI22_X1 U2383 ( .A1(n2135), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[12][10] ), .B2(n2134), .ZN(n2136) );
  INV_X1 U2384 ( .A(n2136), .ZN(n1004) );
  NOR2_X1 U2385 ( .A1(n2247), .A2(n2137), .ZN(n2148) );
  INV_X1 U2386 ( .A(n2148), .ZN(n2149) );
  OAI22_X1 U2387 ( .A1(n2149), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[13][0] ), .B2(n2148), .ZN(n2138) );
  INV_X1 U2388 ( .A(n2138), .ZN(n1003) );
  OAI22_X1 U2389 ( .A1(n2149), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[13][1] ), .B2(n2148), .ZN(n2139) );
  INV_X1 U2390 ( .A(n2139), .ZN(n1002) );
  OAI22_X1 U2391 ( .A1(n2149), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[13][2] ), .B2(n2148), .ZN(n2140) );
  INV_X1 U2392 ( .A(n2140), .ZN(n1001) );
  OAI22_X1 U2393 ( .A1(n2149), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[13][3] ), .B2(n2148), .ZN(n2141) );
  INV_X1 U2394 ( .A(n2141), .ZN(n1000) );
  OAI22_X1 U2395 ( .A1(n2149), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[13][4] ), .B2(n2148), .ZN(n2142) );
  INV_X1 U2396 ( .A(n2142), .ZN(n999) );
  OAI22_X1 U2397 ( .A1(n2149), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[13][5] ), .B2(n2148), .ZN(n2143) );
  INV_X1 U2398 ( .A(n2143), .ZN(n998) );
  OAI22_X1 U2399 ( .A1(n2149), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[13][6] ), .B2(n2148), .ZN(n2144) );
  INV_X1 U2400 ( .A(n2144), .ZN(n997) );
  OAI22_X1 U2401 ( .A1(n2149), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[13][7] ), .B2(n2148), .ZN(n2145) );
  INV_X1 U2402 ( .A(n2145), .ZN(n996) );
  OAI22_X1 U2403 ( .A1(n2149), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[13][8] ), .B2(n2148), .ZN(n2146) );
  INV_X1 U2404 ( .A(n2146), .ZN(n995) );
  OAI22_X1 U2405 ( .A1(n2149), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[13][9] ), .B2(n2148), .ZN(n2147) );
  INV_X1 U2406 ( .A(n2147), .ZN(n994) );
  OAI22_X1 U2407 ( .A1(n2149), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[13][10] ), .B2(n2148), .ZN(n2150) );
  INV_X1 U2408 ( .A(n2150), .ZN(n993) );
  NAND2_X1 U2409 ( .A1(n2276), .A2(n2151), .ZN(n2163) );
  OAI22_X1 U2410 ( .A1(n2163), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[14][0] ), .B2(n2162), .ZN(n2152) );
  INV_X1 U2411 ( .A(n2152), .ZN(n992) );
  OAI22_X1 U2412 ( .A1(n2163), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[14][1] ), .B2(n2162), .ZN(n2153) );
  INV_X1 U2413 ( .A(n2153), .ZN(n991) );
  OAI22_X1 U2414 ( .A1(n2163), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[14][2] ), .B2(n2162), .ZN(n2154) );
  INV_X1 U2415 ( .A(n2154), .ZN(n990) );
  OAI22_X1 U2416 ( .A1(n2163), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[14][3] ), .B2(n2162), .ZN(n2155) );
  INV_X1 U2417 ( .A(n2155), .ZN(n989) );
  OAI22_X1 U2418 ( .A1(n2163), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[14][4] ), .B2(n2162), .ZN(n2156) );
  INV_X1 U2419 ( .A(n2156), .ZN(n988) );
  OAI22_X1 U2420 ( .A1(n2163), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[14][5] ), .B2(n2162), .ZN(n2157) );
  INV_X1 U2421 ( .A(n2157), .ZN(n987) );
  OAI22_X1 U2422 ( .A1(n2163), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[14][6] ), .B2(n2162), .ZN(n2158) );
  INV_X1 U2423 ( .A(n2158), .ZN(n986) );
  OAI22_X1 U2424 ( .A1(n2163), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[14][7] ), .B2(n2162), .ZN(n2159) );
  INV_X1 U2425 ( .A(n2159), .ZN(n985) );
  OAI22_X1 U2426 ( .A1(n2163), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[14][8] ), .B2(n2162), .ZN(n2160) );
  INV_X1 U2427 ( .A(n2160), .ZN(n984) );
  OAI22_X1 U2428 ( .A1(n2163), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[14][9] ), .B2(n2162), .ZN(n2161) );
  INV_X1 U2429 ( .A(n2161), .ZN(n983) );
  OAI22_X1 U2430 ( .A1(n2163), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[14][10] ), .B2(n2162), .ZN(n2164) );
  INV_X1 U2431 ( .A(n2164), .ZN(n982) );
  NOR2_X1 U2432 ( .A1(n2166), .A2(n2165), .ZN(n2177) );
  INV_X1 U2433 ( .A(n2177), .ZN(n2178) );
  OAI22_X1 U2434 ( .A1(n2178), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[15][0] ), .B2(n2177), .ZN(n2167) );
  INV_X1 U2435 ( .A(n2167), .ZN(n981) );
  OAI22_X1 U2436 ( .A1(n2178), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[15][1] ), .B2(n2177), .ZN(n2168) );
  INV_X1 U2437 ( .A(n2168), .ZN(n980) );
  OAI22_X1 U2438 ( .A1(n2178), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[15][2] ), .B2(n2177), .ZN(n2169) );
  INV_X1 U2439 ( .A(n2169), .ZN(n979) );
  OAI22_X1 U2440 ( .A1(n2178), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[15][3] ), .B2(n2177), .ZN(n2170) );
  INV_X1 U2441 ( .A(n2170), .ZN(n978) );
  OAI22_X1 U2442 ( .A1(n2178), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[15][4] ), .B2(n2177), .ZN(n2171) );
  INV_X1 U2443 ( .A(n2171), .ZN(n977) );
  OAI22_X1 U2444 ( .A1(n2178), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[15][5] ), .B2(n2177), .ZN(n2172) );
  INV_X1 U2445 ( .A(n2172), .ZN(n976) );
  OAI22_X1 U2446 ( .A1(n2178), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[15][6] ), .B2(n2177), .ZN(n2173) );
  INV_X1 U2447 ( .A(n2173), .ZN(n975) );
  OAI22_X1 U2448 ( .A1(n2178), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[15][7] ), .B2(n2177), .ZN(n2174) );
  INV_X1 U2449 ( .A(n2174), .ZN(n974) );
  OAI22_X1 U2450 ( .A1(n2178), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[15][8] ), .B2(n2177), .ZN(n2175) );
  INV_X1 U2451 ( .A(n2175), .ZN(n973) );
  OAI22_X1 U2452 ( .A1(n2178), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[15][9] ), .B2(n2177), .ZN(n2176) );
  INV_X1 U2453 ( .A(n2176), .ZN(n972) );
  OAI22_X1 U2454 ( .A1(n2178), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[15][10] ), .B2(n2177), .ZN(n2179) );
  INV_X1 U2455 ( .A(n2179), .ZN(n971) );
  NAND2_X1 U2456 ( .A1(n2276), .A2(n2180), .ZN(n2246) );
  NOR2_X1 U2457 ( .A1(n2290), .A2(n2246), .ZN(n2191) );
  INV_X1 U2458 ( .A(n2191), .ZN(n2192) );
  OAI22_X1 U2459 ( .A1(n2192), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[16][0] ), .B2(n2191), .ZN(n2181) );
  INV_X1 U2460 ( .A(n2181), .ZN(n970) );
  OAI22_X1 U2461 ( .A1(n2192), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[16][1] ), .B2(n2191), .ZN(n2182) );
  INV_X1 U2462 ( .A(n2182), .ZN(n969) );
  OAI22_X1 U2463 ( .A1(n2192), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[16][2] ), .B2(n2191), .ZN(n2183) );
  INV_X1 U2464 ( .A(n2183), .ZN(n968) );
  OAI22_X1 U2465 ( .A1(n2192), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[16][3] ), .B2(n2191), .ZN(n2184) );
  INV_X1 U2466 ( .A(n2184), .ZN(n967) );
  OAI22_X1 U2467 ( .A1(n2192), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[16][4] ), .B2(n2191), .ZN(n2185) );
  INV_X1 U2468 ( .A(n2185), .ZN(n966) );
  OAI22_X1 U2469 ( .A1(n2192), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[16][5] ), .B2(n2191), .ZN(n2186) );
  INV_X1 U2470 ( .A(n2186), .ZN(n965) );
  OAI22_X1 U2471 ( .A1(n2192), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[16][6] ), .B2(n2191), .ZN(n2187) );
  INV_X1 U2472 ( .A(n2187), .ZN(n964) );
  OAI22_X1 U2473 ( .A1(n2192), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[16][7] ), .B2(n2191), .ZN(n2188) );
  INV_X1 U2474 ( .A(n2188), .ZN(n963) );
  OAI22_X1 U2475 ( .A1(n2192), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[16][8] ), .B2(n2191), .ZN(n2189) );
  INV_X1 U2476 ( .A(n2189), .ZN(n962) );
  OAI22_X1 U2477 ( .A1(n2192), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[16][9] ), .B2(n2191), .ZN(n2190) );
  INV_X1 U2478 ( .A(n2190), .ZN(n961) );
  OAI22_X1 U2479 ( .A1(n2192), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[16][10] ), .B2(n2191), .ZN(n2193) );
  INV_X1 U2480 ( .A(n2193), .ZN(n960) );
  NOR2_X1 U2481 ( .A1(n2304), .A2(n2246), .ZN(n2204) );
  INV_X1 U2482 ( .A(n2204), .ZN(n2205) );
  OAI22_X1 U2483 ( .A1(n2205), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[17][0] ), .B2(n2204), .ZN(n2194) );
  INV_X1 U2484 ( .A(n2194), .ZN(n959) );
  OAI22_X1 U2485 ( .A1(n2205), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[17][1] ), .B2(n2204), .ZN(n2195) );
  INV_X1 U2486 ( .A(n2195), .ZN(n958) );
  OAI22_X1 U2487 ( .A1(n2205), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[17][2] ), .B2(n2204), .ZN(n2196) );
  INV_X1 U2488 ( .A(n2196), .ZN(n957) );
  OAI22_X1 U2489 ( .A1(n2205), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[17][3] ), .B2(n2204), .ZN(n2197) );
  INV_X1 U2490 ( .A(n2197), .ZN(n956) );
  OAI22_X1 U2491 ( .A1(n2205), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[17][4] ), .B2(n2204), .ZN(n2198) );
  INV_X1 U2492 ( .A(n2198), .ZN(n955) );
  OAI22_X1 U2493 ( .A1(n2205), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[17][5] ), .B2(n2204), .ZN(n2199) );
  INV_X1 U2494 ( .A(n2199), .ZN(n954) );
  OAI22_X1 U2495 ( .A1(n2205), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[17][6] ), .B2(n2204), .ZN(n2200) );
  INV_X1 U2496 ( .A(n2200), .ZN(n953) );
  OAI22_X1 U2497 ( .A1(n2205), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[17][7] ), .B2(n2204), .ZN(n2201) );
  INV_X1 U2498 ( .A(n2201), .ZN(n952) );
  OAI22_X1 U2499 ( .A1(n2205), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[17][8] ), .B2(n2204), .ZN(n2202) );
  INV_X1 U2500 ( .A(n2202), .ZN(n951) );
  OAI22_X1 U2501 ( .A1(n2205), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[17][9] ), .B2(n2204), .ZN(n2203) );
  INV_X1 U2502 ( .A(n2203), .ZN(n950) );
  OAI22_X1 U2503 ( .A1(n2205), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[17][10] ), .B2(n2204), .ZN(n2206) );
  INV_X1 U2504 ( .A(n2206), .ZN(n949) );
  NOR2_X1 U2505 ( .A1(n2318), .A2(n2246), .ZN(n2217) );
  INV_X1 U2506 ( .A(n2217), .ZN(n2218) );
  OAI22_X1 U2507 ( .A1(n2218), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[18][0] ), .B2(n2217), .ZN(n2207) );
  INV_X1 U2508 ( .A(n2207), .ZN(n948) );
  OAI22_X1 U2509 ( .A1(n2218), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[18][1] ), .B2(n2217), .ZN(n2208) );
  INV_X1 U2510 ( .A(n2208), .ZN(n947) );
  OAI22_X1 U2511 ( .A1(n2218), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[18][2] ), .B2(n2217), .ZN(n2209) );
  INV_X1 U2512 ( .A(n2209), .ZN(n946) );
  OAI22_X1 U2513 ( .A1(n2218), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[18][3] ), .B2(n2217), .ZN(n2210) );
  INV_X1 U2514 ( .A(n2210), .ZN(n945) );
  OAI22_X1 U2515 ( .A1(n2218), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[18][4] ), .B2(n2217), .ZN(n2211) );
  INV_X1 U2516 ( .A(n2211), .ZN(n944) );
  OAI22_X1 U2517 ( .A1(n2218), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[18][5] ), .B2(n2217), .ZN(n2212) );
  INV_X1 U2518 ( .A(n2212), .ZN(n943) );
  OAI22_X1 U2519 ( .A1(n2218), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[18][6] ), .B2(n2217), .ZN(n2213) );
  INV_X1 U2520 ( .A(n2213), .ZN(n942) );
  OAI22_X1 U2521 ( .A1(n2218), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[18][7] ), .B2(n2217), .ZN(n2214) );
  INV_X1 U2522 ( .A(n2214), .ZN(n941) );
  OAI22_X1 U2523 ( .A1(n2218), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[18][8] ), .B2(n2217), .ZN(n2215) );
  INV_X1 U2524 ( .A(n2215), .ZN(n940) );
  OAI22_X1 U2525 ( .A1(n2218), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[18][9] ), .B2(n2217), .ZN(n2216) );
  INV_X1 U2526 ( .A(n2216), .ZN(n939) );
  OAI22_X1 U2527 ( .A1(n2218), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[18][10] ), .B2(n2217), .ZN(n2219) );
  INV_X1 U2528 ( .A(n2219), .ZN(n938) );
  NOR2_X1 U2529 ( .A1(n2332), .A2(n2246), .ZN(n2230) );
  INV_X1 U2530 ( .A(n2230), .ZN(n2231) );
  OAI22_X1 U2531 ( .A1(n2231), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[19][0] ), .B2(n2230), .ZN(n2220) );
  INV_X1 U2532 ( .A(n2220), .ZN(n937) );
  OAI22_X1 U2533 ( .A1(n2231), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[19][1] ), .B2(n2230), .ZN(n2221) );
  INV_X1 U2534 ( .A(n2221), .ZN(n936) );
  OAI22_X1 U2535 ( .A1(n2231), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[19][2] ), .B2(n2230), .ZN(n2222) );
  INV_X1 U2536 ( .A(n2222), .ZN(n935) );
  OAI22_X1 U2537 ( .A1(n2231), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[19][3] ), .B2(n2230), .ZN(n2223) );
  INV_X1 U2538 ( .A(n2223), .ZN(n934) );
  OAI22_X1 U2539 ( .A1(n2231), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[19][4] ), .B2(n2230), .ZN(n2224) );
  INV_X1 U2540 ( .A(n2224), .ZN(n933) );
  OAI22_X1 U2541 ( .A1(n2231), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[19][5] ), .B2(n2230), .ZN(n2225) );
  INV_X1 U2542 ( .A(n2225), .ZN(n932) );
  OAI22_X1 U2543 ( .A1(n2231), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[19][6] ), .B2(n2230), .ZN(n2226) );
  INV_X1 U2544 ( .A(n2226), .ZN(n931) );
  OAI22_X1 U2545 ( .A1(n2231), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[19][7] ), .B2(n2230), .ZN(n2227) );
  INV_X1 U2546 ( .A(n2227), .ZN(n930) );
  OAI22_X1 U2547 ( .A1(n2231), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[19][8] ), .B2(n2230), .ZN(n2228) );
  INV_X1 U2548 ( .A(n2228), .ZN(n929) );
  OAI22_X1 U2549 ( .A1(n2231), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[19][9] ), .B2(n2230), .ZN(n2229) );
  INV_X1 U2550 ( .A(n2229), .ZN(n928) );
  OAI22_X1 U2551 ( .A1(n2231), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[19][10] ), .B2(n2230), .ZN(n2232) );
  INV_X1 U2552 ( .A(n2232), .ZN(n927) );
  NOR2_X1 U2553 ( .A1(n2346), .A2(n2246), .ZN(n2243) );
  INV_X1 U2554 ( .A(n2243), .ZN(n2244) );
  OAI22_X1 U2555 ( .A1(n2244), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[20][0] ), .B2(n2243), .ZN(n2233) );
  INV_X1 U2556 ( .A(n2233), .ZN(n926) );
  OAI22_X1 U2557 ( .A1(n2244), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[20][1] ), .B2(n2243), .ZN(n2234) );
  INV_X1 U2558 ( .A(n2234), .ZN(n925) );
  OAI22_X1 U2559 ( .A1(n2244), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[20][2] ), .B2(n2243), .ZN(n2235) );
  INV_X1 U2560 ( .A(n2235), .ZN(n924) );
  OAI22_X1 U2561 ( .A1(n2244), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[20][3] ), .B2(n2243), .ZN(n2236) );
  INV_X1 U2562 ( .A(n2236), .ZN(n923) );
  OAI22_X1 U2563 ( .A1(n2244), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[20][4] ), .B2(n2243), .ZN(n2237) );
  INV_X1 U2564 ( .A(n2237), .ZN(n922) );
  OAI22_X1 U2565 ( .A1(n2244), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[20][5] ), .B2(n2243), .ZN(n2238) );
  INV_X1 U2566 ( .A(n2238), .ZN(n921) );
  OAI22_X1 U2567 ( .A1(n2244), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[20][6] ), .B2(n2243), .ZN(n2239) );
  INV_X1 U2568 ( .A(n2239), .ZN(n920) );
  OAI22_X1 U2569 ( .A1(n2244), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[20][7] ), .B2(n2243), .ZN(n2240) );
  INV_X1 U2570 ( .A(n2240), .ZN(n919) );
  OAI22_X1 U2571 ( .A1(n2244), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[20][8] ), .B2(n2243), .ZN(n2241) );
  INV_X1 U2572 ( .A(n2241), .ZN(n918) );
  OAI22_X1 U2573 ( .A1(n2244), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[20][9] ), .B2(n2243), .ZN(n2242) );
  INV_X1 U2574 ( .A(n2242), .ZN(n917) );
  OAI22_X1 U2575 ( .A1(n2244), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[20][10] ), .B2(n2243), .ZN(n2245) );
  INV_X1 U2576 ( .A(n2245), .ZN(n916) );
  NOR2_X1 U2577 ( .A1(n2247), .A2(n2246), .ZN(n2258) );
  INV_X1 U2578 ( .A(n2258), .ZN(n2259) );
  OAI22_X1 U2579 ( .A1(n2259), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[21][0] ), .B2(n2258), .ZN(n2248) );
  INV_X1 U2580 ( .A(n2248), .ZN(n915) );
  OAI22_X1 U2581 ( .A1(n2259), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[21][1] ), .B2(n2258), .ZN(n2249) );
  INV_X1 U2582 ( .A(n2249), .ZN(n914) );
  OAI22_X1 U2583 ( .A1(n2259), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[21][2] ), .B2(n2258), .ZN(n2250) );
  INV_X1 U2584 ( .A(n2250), .ZN(n913) );
  OAI22_X1 U2585 ( .A1(n2259), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[21][3] ), .B2(n2258), .ZN(n2251) );
  INV_X1 U2586 ( .A(n2251), .ZN(n912) );
  OAI22_X1 U2587 ( .A1(n2259), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[21][4] ), .B2(n2258), .ZN(n2252) );
  INV_X1 U2588 ( .A(n2252), .ZN(n911) );
  OAI22_X1 U2589 ( .A1(n2259), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[21][5] ), .B2(n2258), .ZN(n2253) );
  INV_X1 U2590 ( .A(n2253), .ZN(n910) );
  OAI22_X1 U2591 ( .A1(n2259), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[21][6] ), .B2(n2258), .ZN(n2254) );
  INV_X1 U2592 ( .A(n2254), .ZN(n909) );
  OAI22_X1 U2593 ( .A1(n2259), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[21][7] ), .B2(n2258), .ZN(n2255) );
  INV_X1 U2594 ( .A(n2255), .ZN(n908) );
  OAI22_X1 U2595 ( .A1(n2259), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[21][8] ), .B2(n2258), .ZN(n2256) );
  INV_X1 U2596 ( .A(n2256), .ZN(n907) );
  OAI22_X1 U2597 ( .A1(n2259), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[21][9] ), .B2(n2258), .ZN(n2257) );
  INV_X1 U2598 ( .A(n2257), .ZN(n906) );
  OAI22_X1 U2599 ( .A1(n2259), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[21][10] ), .B2(n2258), .ZN(n2260) );
  INV_X1 U2600 ( .A(n2260), .ZN(n905) );
  NAND2_X1 U2601 ( .A1(n2276), .A2(n2261), .ZN(n2273) );
  OAI22_X1 U2602 ( .A1(n2273), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[22][0] ), .B2(n2272), .ZN(n2262) );
  INV_X1 U2603 ( .A(n2262), .ZN(n904) );
  OAI22_X1 U2604 ( .A1(n2273), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[22][1] ), .B2(n2272), .ZN(n2263) );
  INV_X1 U2605 ( .A(n2263), .ZN(n903) );
  OAI22_X1 U2606 ( .A1(n2273), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[22][2] ), .B2(n2272), .ZN(n2264) );
  INV_X1 U2607 ( .A(n2264), .ZN(n902) );
  OAI22_X1 U2608 ( .A1(n2273), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[22][3] ), .B2(n2272), .ZN(n2265) );
  INV_X1 U2609 ( .A(n2265), .ZN(n901) );
  OAI22_X1 U2610 ( .A1(n2273), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[22][4] ), .B2(n2272), .ZN(n2266) );
  INV_X1 U2611 ( .A(n2266), .ZN(n900) );
  OAI22_X1 U2612 ( .A1(n2273), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[22][5] ), .B2(n2272), .ZN(n2267) );
  INV_X1 U2613 ( .A(n2267), .ZN(n899) );
  OAI22_X1 U2614 ( .A1(n2273), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[22][6] ), .B2(n2272), .ZN(n2268) );
  INV_X1 U2615 ( .A(n2268), .ZN(n898) );
  OAI22_X1 U2616 ( .A1(n2273), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[22][7] ), .B2(n2272), .ZN(n2269) );
  INV_X1 U2617 ( .A(n2269), .ZN(n897) );
  OAI22_X1 U2618 ( .A1(n2273), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[22][8] ), .B2(n2272), .ZN(n2270) );
  INV_X1 U2619 ( .A(n2270), .ZN(n896) );
  OAI22_X1 U2620 ( .A1(n2273), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[22][9] ), .B2(n2272), .ZN(n2271) );
  INV_X1 U2621 ( .A(n2271), .ZN(n895) );
  OAI22_X1 U2622 ( .A1(n2273), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[22][10] ), .B2(n2272), .ZN(n2274) );
  INV_X1 U2623 ( .A(n2274), .ZN(n894) );
  NAND2_X1 U2624 ( .A1(n2276), .A2(n2275), .ZN(n2288) );
  INV_X1 U2625 ( .A(n2288), .ZN(n2287) );
  OAI22_X1 U2626 ( .A1(n2288), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[23][0] ), .B2(n2287), .ZN(n2277) );
  INV_X1 U2627 ( .A(n2277), .ZN(n893) );
  OAI22_X1 U2628 ( .A1(n2288), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[23][1] ), .B2(n2287), .ZN(n2278) );
  INV_X1 U2629 ( .A(n2278), .ZN(n892) );
  OAI22_X1 U2630 ( .A1(n2288), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[23][2] ), .B2(n2287), .ZN(n2279) );
  INV_X1 U2631 ( .A(n2279), .ZN(n891) );
  OAI22_X1 U2632 ( .A1(n2288), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[23][3] ), .B2(n2287), .ZN(n2280) );
  INV_X1 U2633 ( .A(n2280), .ZN(n890) );
  OAI22_X1 U2634 ( .A1(n2288), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[23][4] ), .B2(n2287), .ZN(n2281) );
  INV_X1 U2635 ( .A(n2281), .ZN(n889) );
  OAI22_X1 U2636 ( .A1(n2288), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[23][5] ), .B2(n2287), .ZN(n2282) );
  INV_X1 U2637 ( .A(n2282), .ZN(n888) );
  OAI22_X1 U2638 ( .A1(n2288), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[23][6] ), .B2(n2287), .ZN(n2283) );
  INV_X1 U2639 ( .A(n2283), .ZN(n887) );
  OAI22_X1 U2640 ( .A1(n2288), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[23][7] ), .B2(n2287), .ZN(n2284) );
  INV_X1 U2641 ( .A(n2284), .ZN(n886) );
  OAI22_X1 U2642 ( .A1(n2288), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[23][8] ), .B2(n2287), .ZN(n2285) );
  INV_X1 U2643 ( .A(n2285), .ZN(n885) );
  OAI22_X1 U2644 ( .A1(n2288), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[23][9] ), .B2(n2287), .ZN(n2286) );
  INV_X1 U2645 ( .A(n2286), .ZN(n884) );
  OAI22_X1 U2646 ( .A1(n2288), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[23][10] ), .B2(n2287), .ZN(n2289) );
  INV_X1 U2647 ( .A(n2289), .ZN(n883) );
  NOR2_X1 U2648 ( .A1(n2347), .A2(n2290), .ZN(n2301) );
  INV_X1 U2649 ( .A(n2301), .ZN(n2302) );
  OAI22_X1 U2650 ( .A1(n2302), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[24][0] ), .B2(n2301), .ZN(n2291) );
  INV_X1 U2651 ( .A(n2291), .ZN(n882) );
  OAI22_X1 U2652 ( .A1(n2302), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[24][1] ), .B2(n2301), .ZN(n2292) );
  INV_X1 U2653 ( .A(n2292), .ZN(n881) );
  OAI22_X1 U2654 ( .A1(n2302), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[24][2] ), .B2(n2301), .ZN(n2293) );
  INV_X1 U2655 ( .A(n2293), .ZN(n880) );
  OAI22_X1 U2656 ( .A1(n2302), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[24][3] ), .B2(n2301), .ZN(n2294) );
  INV_X1 U2657 ( .A(n2294), .ZN(n879) );
  OAI22_X1 U2658 ( .A1(n2302), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[24][4] ), .B2(n2301), .ZN(n2295) );
  INV_X1 U2659 ( .A(n2295), .ZN(n878) );
  OAI22_X1 U2660 ( .A1(n2302), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[24][5] ), .B2(n2301), .ZN(n2296) );
  INV_X1 U2661 ( .A(n2296), .ZN(n877) );
  OAI22_X1 U2662 ( .A1(n2302), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[24][6] ), .B2(n2301), .ZN(n2297) );
  INV_X1 U2663 ( .A(n2297), .ZN(n876) );
  OAI22_X1 U2664 ( .A1(n2302), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[24][7] ), .B2(n2301), .ZN(n2298) );
  INV_X1 U2665 ( .A(n2298), .ZN(n875) );
  OAI22_X1 U2666 ( .A1(n2302), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[24][8] ), .B2(n2301), .ZN(n2299) );
  INV_X1 U2667 ( .A(n2299), .ZN(n874) );
  OAI22_X1 U2668 ( .A1(n2302), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[24][9] ), .B2(n2301), .ZN(n2300) );
  INV_X1 U2669 ( .A(n2300), .ZN(n873) );
  OAI22_X1 U2670 ( .A1(n2302), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[24][10] ), .B2(n2301), .ZN(n2303) );
  INV_X1 U2671 ( .A(n2303), .ZN(n872) );
  NOR2_X1 U2672 ( .A1(n2347), .A2(n2304), .ZN(n2315) );
  INV_X1 U2673 ( .A(n2315), .ZN(n2316) );
  OAI22_X1 U2674 ( .A1(n2316), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[25][0] ), .B2(n2315), .ZN(n2305) );
  INV_X1 U2675 ( .A(n2305), .ZN(n871) );
  OAI22_X1 U2676 ( .A1(n2316), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[25][1] ), .B2(n2315), .ZN(n2306) );
  INV_X1 U2677 ( .A(n2306), .ZN(n870) );
  OAI22_X1 U2678 ( .A1(n2316), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[25][2] ), .B2(n2315), .ZN(n2307) );
  INV_X1 U2679 ( .A(n2307), .ZN(n869) );
  OAI22_X1 U2680 ( .A1(n2316), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[25][3] ), .B2(n2315), .ZN(n2308) );
  INV_X1 U2681 ( .A(n2308), .ZN(n868) );
  OAI22_X1 U2682 ( .A1(n2316), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[25][4] ), .B2(n2315), .ZN(n2309) );
  INV_X1 U2683 ( .A(n2309), .ZN(n867) );
  OAI22_X1 U2684 ( .A1(n2316), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[25][5] ), .B2(n2315), .ZN(n2310) );
  INV_X1 U2685 ( .A(n2310), .ZN(n866) );
  OAI22_X1 U2686 ( .A1(n2316), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[25][6] ), .B2(n2315), .ZN(n2311) );
  INV_X1 U2687 ( .A(n2311), .ZN(n865) );
  OAI22_X1 U2688 ( .A1(n2316), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[25][7] ), .B2(n2315), .ZN(n2312) );
  INV_X1 U2689 ( .A(n2312), .ZN(n864) );
  OAI22_X1 U2690 ( .A1(n2316), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[25][8] ), .B2(n2315), .ZN(n2313) );
  INV_X1 U2691 ( .A(n2313), .ZN(n863) );
  OAI22_X1 U2692 ( .A1(n2316), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[25][9] ), .B2(n2315), .ZN(n2314) );
  INV_X1 U2693 ( .A(n2314), .ZN(n862) );
  OAI22_X1 U2694 ( .A1(n2316), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[25][10] ), .B2(n2315), .ZN(n2317) );
  INV_X1 U2695 ( .A(n2317), .ZN(n861) );
  NOR2_X1 U2696 ( .A1(n2347), .A2(n2318), .ZN(n2329) );
  INV_X1 U2697 ( .A(n2329), .ZN(n2330) );
  OAI22_X1 U2698 ( .A1(n2330), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[26][0] ), .B2(n2329), .ZN(n2319) );
  INV_X1 U2699 ( .A(n2319), .ZN(n860) );
  OAI22_X1 U2700 ( .A1(n2330), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[26][1] ), .B2(n2329), .ZN(n2320) );
  INV_X1 U2701 ( .A(n2320), .ZN(n859) );
  OAI22_X1 U2702 ( .A1(n2330), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[26][2] ), .B2(n2329), .ZN(n2321) );
  INV_X1 U2703 ( .A(n2321), .ZN(n858) );
  OAI22_X1 U2704 ( .A1(n2330), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[26][3] ), .B2(n2329), .ZN(n2322) );
  INV_X1 U2705 ( .A(n2322), .ZN(n857) );
  OAI22_X1 U2706 ( .A1(n2330), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[26][4] ), .B2(n2329), .ZN(n2323) );
  INV_X1 U2707 ( .A(n2323), .ZN(n856) );
  OAI22_X1 U2708 ( .A1(n2330), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[26][5] ), .B2(n2329), .ZN(n2324) );
  INV_X1 U2709 ( .A(n2324), .ZN(n855) );
  OAI22_X1 U2710 ( .A1(n2330), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[26][6] ), .B2(n2329), .ZN(n2325) );
  INV_X1 U2711 ( .A(n2325), .ZN(n854) );
  OAI22_X1 U2712 ( .A1(n2330), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[26][7] ), .B2(n2329), .ZN(n2326) );
  INV_X1 U2713 ( .A(n2326), .ZN(n853) );
  OAI22_X1 U2714 ( .A1(n2330), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[26][8] ), .B2(n2329), .ZN(n2327) );
  INV_X1 U2715 ( .A(n2327), .ZN(n852) );
  OAI22_X1 U2716 ( .A1(n2330), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[26][9] ), .B2(n2329), .ZN(n2328) );
  INV_X1 U2717 ( .A(n2328), .ZN(n851) );
  OAI22_X1 U2718 ( .A1(n2330), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[26][10] ), .B2(n2329), .ZN(n2331) );
  INV_X1 U2719 ( .A(n2331), .ZN(n850) );
  NOR2_X1 U2720 ( .A1(n2347), .A2(n2332), .ZN(n2343) );
  INV_X1 U2721 ( .A(n2343), .ZN(n2344) );
  OAI22_X1 U2722 ( .A1(n2344), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[27][0] ), .B2(n2343), .ZN(n2333) );
  INV_X1 U2723 ( .A(n2333), .ZN(n849) );
  OAI22_X1 U2724 ( .A1(n2344), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[27][1] ), .B2(n2343), .ZN(n2334) );
  INV_X1 U2725 ( .A(n2334), .ZN(n848) );
  OAI22_X1 U2726 ( .A1(n2344), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[27][2] ), .B2(n2343), .ZN(n2335) );
  INV_X1 U2727 ( .A(n2335), .ZN(n847) );
  OAI22_X1 U2728 ( .A1(n2344), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[27][3] ), .B2(n2343), .ZN(n2336) );
  INV_X1 U2729 ( .A(n2336), .ZN(n846) );
  OAI22_X1 U2730 ( .A1(n2344), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[27][4] ), .B2(n2343), .ZN(n2337) );
  INV_X1 U2731 ( .A(n2337), .ZN(n845) );
  OAI22_X1 U2732 ( .A1(n2344), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[27][5] ), .B2(n2343), .ZN(n2338) );
  INV_X1 U2733 ( .A(n2338), .ZN(n844) );
  OAI22_X1 U2734 ( .A1(n2344), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[27][6] ), .B2(n2343), .ZN(n2339) );
  INV_X1 U2735 ( .A(n2339), .ZN(n843) );
  OAI22_X1 U2736 ( .A1(n2344), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[27][7] ), .B2(n2343), .ZN(n2340) );
  INV_X1 U2737 ( .A(n2340), .ZN(n842) );
  OAI22_X1 U2738 ( .A1(n2344), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[27][8] ), .B2(n2343), .ZN(n2341) );
  INV_X1 U2739 ( .A(n2341), .ZN(n841) );
  OAI22_X1 U2740 ( .A1(n2344), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[27][9] ), .B2(n2343), .ZN(n2342) );
  INV_X1 U2741 ( .A(n2342), .ZN(n840) );
  OAI22_X1 U2742 ( .A1(n2344), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[27][10] ), .B2(n2343), .ZN(n2345) );
  INV_X1 U2743 ( .A(n2345), .ZN(n839) );
  NOR2_X1 U2744 ( .A1(n2347), .A2(n2346), .ZN(n2358) );
  INV_X1 U2745 ( .A(n2358), .ZN(n2359) );
  OAI22_X1 U2746 ( .A1(n2359), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[28][0] ), .B2(n2358), .ZN(n2348) );
  INV_X1 U2747 ( .A(n2348), .ZN(n838) );
  OAI22_X1 U2748 ( .A1(n2359), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[28][1] ), .B2(n2358), .ZN(n2349) );
  INV_X1 U2749 ( .A(n2349), .ZN(n837) );
  OAI22_X1 U2750 ( .A1(n2359), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[28][2] ), .B2(n2358), .ZN(n2350) );
  INV_X1 U2751 ( .A(n2350), .ZN(n836) );
  OAI22_X1 U2752 ( .A1(n2359), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[28][3] ), .B2(n2358), .ZN(n2351) );
  INV_X1 U2753 ( .A(n2351), .ZN(n835) );
  OAI22_X1 U2754 ( .A1(n2359), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[28][4] ), .B2(n2358), .ZN(n2352) );
  INV_X1 U2755 ( .A(n2352), .ZN(n834) );
  OAI22_X1 U2756 ( .A1(n2359), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[28][5] ), .B2(n2358), .ZN(n2353) );
  INV_X1 U2757 ( .A(n2353), .ZN(n833) );
  OAI22_X1 U2758 ( .A1(n2359), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[28][6] ), .B2(n2358), .ZN(n2354) );
  INV_X1 U2759 ( .A(n2354), .ZN(n832) );
  OAI22_X1 U2760 ( .A1(n2359), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[28][7] ), .B2(n2358), .ZN(n2355) );
  INV_X1 U2761 ( .A(n2355), .ZN(n831) );
  OAI22_X1 U2762 ( .A1(n2359), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[28][8] ), .B2(n2358), .ZN(n2356) );
  INV_X1 U2763 ( .A(n2356), .ZN(n830) );
  OAI22_X1 U2764 ( .A1(n2359), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[28][9] ), .B2(n2358), .ZN(n2357) );
  INV_X1 U2765 ( .A(n2357), .ZN(n829) );
  OAI22_X1 U2766 ( .A1(n2359), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[28][10] ), .B2(n2358), .ZN(n2360) );
  INV_X1 U2767 ( .A(n2360), .ZN(n828) );
  INV_X1 U2768 ( .A(n2371), .ZN(n2372) );
  OAI22_X1 U2769 ( .A1(n2372), .A2(s_data_in_x[0]), .B1(\xmem_inst/mem[29][0] ), .B2(n2371), .ZN(n2361) );
  INV_X1 U2770 ( .A(n2361), .ZN(n827) );
  OAI22_X1 U2771 ( .A1(n2372), .A2(s_data_in_x[1]), .B1(\xmem_inst/mem[29][1] ), .B2(n2371), .ZN(n2362) );
  INV_X1 U2772 ( .A(n2362), .ZN(n826) );
  OAI22_X1 U2773 ( .A1(n2372), .A2(s_data_in_x[2]), .B1(\xmem_inst/mem[29][2] ), .B2(n2371), .ZN(n2363) );
  INV_X1 U2774 ( .A(n2363), .ZN(n825) );
  OAI22_X1 U2775 ( .A1(n2372), .A2(s_data_in_x[3]), .B1(\xmem_inst/mem[29][3] ), .B2(n2371), .ZN(n2364) );
  INV_X1 U2776 ( .A(n2364), .ZN(n824) );
  OAI22_X1 U2777 ( .A1(n2372), .A2(s_data_in_x[4]), .B1(\xmem_inst/mem[29][4] ), .B2(n2371), .ZN(n2365) );
  INV_X1 U2778 ( .A(n2365), .ZN(n823) );
  OAI22_X1 U2779 ( .A1(n2372), .A2(s_data_in_x[5]), .B1(\xmem_inst/mem[29][5] ), .B2(n2371), .ZN(n2366) );
  INV_X1 U2780 ( .A(n2366), .ZN(n822) );
  OAI22_X1 U2781 ( .A1(n2372), .A2(s_data_in_x[6]), .B1(\xmem_inst/mem[29][6] ), .B2(n2371), .ZN(n2367) );
  INV_X1 U2782 ( .A(n2367), .ZN(n821) );
  OAI22_X1 U2783 ( .A1(n2372), .A2(s_data_in_x[7]), .B1(\xmem_inst/mem[29][7] ), .B2(n2371), .ZN(n2368) );
  INV_X1 U2784 ( .A(n2368), .ZN(n820) );
  OAI22_X1 U2785 ( .A1(n2372), .A2(s_data_in_x[8]), .B1(\xmem_inst/mem[29][8] ), .B2(n2371), .ZN(n2369) );
  INV_X1 U2786 ( .A(n2369), .ZN(n819) );
  OAI22_X1 U2787 ( .A1(n2372), .A2(s_data_in_x[9]), .B1(\xmem_inst/mem[29][9] ), .B2(n2371), .ZN(n2370) );
  INV_X1 U2788 ( .A(n2370), .ZN(n818) );
  OAI22_X1 U2789 ( .A1(n2372), .A2(s_data_in_x[10]), .B1(
        \xmem_inst/mem[29][10] ), .B2(n2371), .ZN(n2373) );
  INV_X1 U2790 ( .A(n2373), .ZN(n817) );
  OAI21_X1 U2791 ( .B1(n2496), .B2(n2375), .A(n2374), .ZN(n816) );
  NAND2_X1 U2792 ( .A1(fmem_addr[1]), .A2(fmem_addr[0]), .ZN(n2376) );
  OAI22_X1 U2793 ( .A1(n2378), .A2(n2489), .B1(n2377), .B2(n2376), .ZN(n814)
         );
  OAI22_X1 U2794 ( .A1(n2490), .A2(n2380), .B1(n2379), .B2(n2503), .ZN(n806)
         );
  NAND2_X1 U2795 ( .A1(m_valid_y), .A2(n2381), .ZN(n2469) );
  INV_X1 U2796 ( .A(n2469), .ZN(n2462) );
  NOR2_X1 U2797 ( .A1(n2483), .A2(n2520), .ZN(n2382) );
  NAND2_X1 U2798 ( .A1(n2382), .A2(\mac_unit_inst/adder_reg [1]), .ZN(n2419)
         );
  OR2_X1 U2799 ( .A1(n2481), .A2(n2517), .ZN(n2418) );
  NAND2_X1 U2800 ( .A1(n2480), .A2(\mac_unit_inst/x_mult_f_reg [2]), .ZN(n2383) );
  AND2_X1 U2801 ( .A1(n2418), .A2(n2383), .ZN(n2384) );
  AND2_X1 U2802 ( .A1(n2419), .A2(n2384), .ZN(n2387) );
  NOR2_X1 U2803 ( .A1(n2483), .A2(n2520), .ZN(n2385) );
  NAND2_X1 U2804 ( .A1(n2385), .A2(\mac_unit_inst/x_mult_f_reg [1]), .ZN(n2420) );
  NOR2_X1 U2805 ( .A1(\mac_unit_inst/x_mult_f_reg [2]), .A2(n2480), .ZN(n2386)
         );
  AOI21_X1 U2806 ( .B1(n2387), .B2(n2420), .A(n2386), .ZN(n2426) );
  NAND2_X1 U2807 ( .A1(n2429), .A2(n1237), .ZN(n2389) );
  NAND2_X1 U2808 ( .A1(\mac_unit_inst/adder_reg [4]), .A2(
        \mac_unit_inst/x_mult_f_reg [4]), .ZN(n2388) );
  NAND2_X1 U2809 ( .A1(n2389), .A2(n2388), .ZN(n2433) );
  INV_X1 U2810 ( .A(n2443), .ZN(n2452) );
  NOR2_X1 U2811 ( .A1(\mac_unit_inst/x_mult_f_reg [6]), .A2(
        \mac_unit_inst/adder_reg [6]), .ZN(n2394) );
  INV_X1 U2812 ( .A(n2394), .ZN(n2442) );
  NAND2_X1 U2813 ( .A1(\mac_unit_inst/adder_reg [6]), .A2(
        \mac_unit_inst/x_mult_f_reg [6]), .ZN(n2390) );
  INV_X1 U2814 ( .A(n2390), .ZN(n2441) );
  NOR2_X1 U2815 ( .A1(n2390), .A2(n1222), .ZN(n2392) );
  AND2_X1 U2816 ( .A1(\mac_unit_inst/adder_reg [7]), .A2(
        \mac_unit_inst/x_mult_f_reg [7]), .ZN(n2391) );
  OR2_X1 U2817 ( .A1(n2392), .A2(n2391), .ZN(n2393) );
  AOI21_X1 U2818 ( .B1(n1223), .B2(n2441), .A(n2393), .ZN(n2450) );
  NAND2_X1 U2819 ( .A1(\mac_unit_inst/adder_reg [9]), .A2(
        \mac_unit_inst/x_mult_f_reg [9]), .ZN(n2396) );
  NAND2_X1 U2820 ( .A1(\mac_unit_inst/adder_reg [8]), .A2(
        \mac_unit_inst/x_mult_f_reg [8]), .ZN(n2457) );
  NOR2_X1 U2821 ( .A1(n2394), .A2(n1222), .ZN(n2395) );
  NOR2_X1 U2822 ( .A1(n1223), .A2(n2395), .ZN(n2451) );
  NAND2_X1 U2823 ( .A1(n2397), .A2(n2396), .ZN(n2398) );
  INV_X1 U2824 ( .A(\mac_unit_inst/x_mult_f_reg [10]), .ZN(n2405) );
  NAND2_X1 U2825 ( .A1(n2411), .A2(n2405), .ZN(n2404) );
  NAND2_X1 U2826 ( .A1(n2411), .A2(n2488), .ZN(n2403) );
  NAND2_X1 U2827 ( .A1(n2405), .A2(n2488), .ZN(n2402) );
  NAND3_X1 U2828 ( .A1(n2404), .A2(n2403), .A3(n2402), .ZN(n2412) );
  XNOR2_X1 U2829 ( .A(n2405), .B(n2488), .ZN(n2410) );
  XNOR2_X1 U2830 ( .A(n2411), .B(n2410), .ZN(n2406) );
  NOR2_X1 U2831 ( .A1(m_valid_y), .A2(n2505), .ZN(n2408) );
  NAND2_X1 U2832 ( .A1(n2408), .A2(n2407), .ZN(n2425) );
  NOR2_X1 U2833 ( .A1(n2467), .A2(n2425), .ZN(n2439) );
  XOR2_X1 U2834 ( .A(\mac_unit_inst/adder_reg [0]), .B(
        \mac_unit_inst/x_mult_f_reg [0]), .Z(n2409) );
  AOI22_X1 U2835 ( .A1(n2462), .A2(\mac_unit_inst/adder_reg [0]), .B1(n2439), 
        .B2(n2409), .ZN(n2413) );
  AND2_X1 U2836 ( .A1(n2412), .A2(n2406), .ZN(n2471) );
  INV_X1 U2837 ( .A(n2425), .ZN(n2468) );
  NAND2_X1 U2838 ( .A1(n2413), .A2(n2465), .ZN(n794) );
  NOR2_X1 U2839 ( .A1(n2467), .A2(n2425), .ZN(n2435) );
  NOR2_X1 U2840 ( .A1(n2483), .A2(n2520), .ZN(n2415) );
  XOR2_X1 U2841 ( .A(\mac_unit_inst/adder_reg [1]), .B(
        \mac_unit_inst/x_mult_f_reg [1]), .Z(n2414) );
  XOR2_X1 U2842 ( .A(n2415), .B(n2414), .Z(n2416) );
  AOI22_X1 U2843 ( .A1(n2462), .A2(\mac_unit_inst/adder_reg [1]), .B1(n2435), 
        .B2(n2416), .ZN(n2417) );
  NAND2_X1 U2844 ( .A1(n2417), .A2(n2465), .ZN(n793) );
  NOR2_X1 U2845 ( .A1(n2467), .A2(n2425), .ZN(n2448) );
  NAND3_X1 U2846 ( .A1(n2420), .A2(n2419), .A3(n2418), .ZN(n2422) );
  XOR2_X1 U2847 ( .A(n2480), .B(\mac_unit_inst/x_mult_f_reg [2]), .Z(n2421) );
  XOR2_X1 U2848 ( .A(n2422), .B(n2421), .Z(n2423) );
  AOI22_X1 U2849 ( .A1(n2462), .A2(n2480), .B1(n2448), .B2(n2423), .ZN(n2424)
         );
  NAND2_X1 U2850 ( .A1(n2424), .A2(n2465), .ZN(n792) );
  NOR2_X1 U2851 ( .A1(n2467), .A2(n2425), .ZN(n2464) );
  FA_X1 U2852 ( .A(\mac_unit_inst/adder_reg [3]), .B(
        \mac_unit_inst/x_mult_f_reg [3]), .CI(n2426), .CO(n2429), .S(n2427) );
  AOI21_X1 U2853 ( .B1(n2464), .B2(n2427), .A(n1226), .ZN(n2428) );
  NAND2_X1 U2854 ( .A1(n2428), .A2(n2465), .ZN(n791) );
  XOR2_X1 U2855 ( .A(\mac_unit_inst/adder_reg [4]), .B(
        \mac_unit_inst/x_mult_f_reg [4]), .Z(n2430) );
  XOR2_X1 U2856 ( .A(n2429), .B(n2430), .Z(n2431) );
  AOI22_X1 U2857 ( .A1(n2462), .A2(\mac_unit_inst/adder_reg [4]), .B1(n2448), 
        .B2(n2431), .ZN(n2432) );
  NAND2_X1 U2858 ( .A1(n2432), .A2(n2465), .ZN(n790) );
  FA_X1 U2859 ( .A(\mac_unit_inst/adder_reg [5]), .B(
        \mac_unit_inst/x_mult_f_reg [5]), .CI(n2433), .CO(n2443), .S(n2434) );
  AOI22_X1 U2860 ( .A1(n2462), .A2(\mac_unit_inst/adder_reg [5]), .B1(n2435), 
        .B2(n2434), .ZN(n2436) );
  NAND2_X1 U2861 ( .A1(n2436), .A2(n2465), .ZN(n789) );
  XOR2_X1 U2862 ( .A(\mac_unit_inst/adder_reg [6]), .B(
        \mac_unit_inst/x_mult_f_reg [6]), .Z(n2437) );
  XOR2_X1 U2863 ( .A(n2443), .B(n2437), .Z(n2438) );
  AOI22_X1 U2864 ( .A1(n2462), .A2(\mac_unit_inst/adder_reg [6]), .B1(n2439), 
        .B2(n2438), .ZN(n2440) );
  NAND2_X1 U2865 ( .A1(n2440), .A2(n2465), .ZN(n788) );
  AOI21_X1 U2866 ( .B1(n2443), .B2(n2442), .A(n2441), .ZN(n2444) );
  INV_X1 U2867 ( .A(n2444), .ZN(n2446) );
  XOR2_X1 U2868 ( .A(\mac_unit_inst/adder_reg [7]), .B(
        \mac_unit_inst/x_mult_f_reg [7]), .Z(n2445) );
  XOR2_X1 U2869 ( .A(n2446), .B(n2445), .Z(n2447) );
  AOI22_X1 U2870 ( .A1(n2462), .A2(\mac_unit_inst/adder_reg [7]), .B1(n2448), 
        .B2(n2447), .ZN(n2449) );
  NAND2_X1 U2871 ( .A1(n2449), .A2(n2465), .ZN(n787) );
  XOR2_X1 U2872 ( .A(\mac_unit_inst/adder_reg [8]), .B(
        \mac_unit_inst/x_mult_f_reg [8]), .Z(n2453) );
  XOR2_X1 U2873 ( .A(n2456), .B(n2453), .Z(n2454) );
  NAND2_X1 U2874 ( .A1(n2455), .A2(n2465), .ZN(n786) );
  NAND3_X1 U2875 ( .A1(n2459), .A2(n2458), .A3(n2457), .ZN(n2461) );
  XOR2_X1 U2876 ( .A(\mac_unit_inst/adder_reg [9]), .B(
        \mac_unit_inst/x_mult_f_reg [9]), .Z(n2460) );
  XOR2_X1 U2877 ( .A(n2461), .B(n2460), .Z(n2463) );
  AOI21_X1 U2878 ( .B1(n2464), .B2(n2463), .A(n1239), .ZN(n2466) );
  NAND2_X1 U2879 ( .A1(n2466), .A2(n2465), .ZN(n785) );
  OAI21_X1 U2880 ( .B1(n2467), .B2(n2406), .A(n2468), .ZN(n2470) );
  OAI22_X1 U2881 ( .A1(n2471), .A2(n2470), .B1(n2488), .B2(n2469), .ZN(n784)
         );
endmodule

